-- Computer_System.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Computer_System is
	port (
		arduino_gpio_export             : inout std_logic_vector(15 downto 0) := (others => '0'); --            arduino_gpio.export
		arduino_reset_n_export          : out   std_logic;                                        --         arduino_reset_n.export
		blinky_export                   : out   std_logic;                                        --                  blinky.export
		expansion_jp1_export            : inout std_logic_vector(31 downto 0) := (others => '0'); --           expansion_jp1.export
		hex3_hex0_export                : out   std_logic_vector(31 downto 0);                    --               hex3_hex0.export
		hex5_hex4_export                : out   std_logic_vector(31 downto 0);                    --               hex5_hex4.export
		iservo_control_0_export         : out   std_logic_vector(15 downto 0);                    --        iservo_control_0.export
		iservo_control_1_export         : out   std_logic_vector(15 downto 0);                    --        iservo_control_1.export
		leds_export                     : out   std_logic_vector(9 downto 0);                     --                    leds.export
		pushbuttons_export              : in    std_logic_vector(1 downto 0)  := (others => '0'); --             pushbuttons.export
		sdram_addr                      : out   std_logic_vector(12 downto 0);                    --                   sdram.addr
		sdram_ba                        : out   std_logic_vector(1 downto 0);                     --                        .ba
		sdram_cas_n                     : out   std_logic;                                        --                        .cas_n
		sdram_cke                       : out   std_logic;                                        --                        .cke
		sdram_cs_n                      : out   std_logic;                                        --                        .cs_n
		sdram_dq                        : inout std_logic_vector(15 downto 0) := (others => '0'); --                        .dq
		sdram_dqm                       : out   std_logic_vector(1 downto 0);                     --                        .dqm
		sdram_ras_n                     : out   std_logic;                                        --                        .ras_n
		sdram_we_n                      : out   std_logic;                                        --                        .we_n
		sdram_clk_clk                   : out   std_logic;                                        --               sdram_clk.clk
		servo_control_0_export          : out   std_logic;                                        --         servo_control_0.export
		servo_control_1_export          : out   std_logic;                                        --         servo_control_1.export
		slider_switches_export          : in    std_logic_vector(9 downto 0)  := (others => '0'); --         slider_switches.export
		system_pll_ref_clk_clk          : in    std_logic                     := '0';             --      system_pll_ref_clk.clk
		system_pll_ref_reset_reset      : in    std_logic                     := '0';             --    system_pll_ref_reset.reset
		video_lt24_controller_0_lcd_on  : out   std_logic;                                        -- video_lt24_controller_0.lcd_on
		video_lt24_controller_0_reset_n : out   std_logic;                                        --                        .reset_n
		video_lt24_controller_0_csx     : out   std_logic;                                        --                        .csx
		video_lt24_controller_0_data    : out   std_logic_vector(15 downto 0);                    --                        .data
		video_lt24_controller_0_rdx     : out   std_logic;                                        --                        .rdx
		video_lt24_controller_0_wrx     : out   std_logic;                                        --                        .wrx
		video_lt24_controller_0_dcx     : out   std_logic;                                        --                        .dcx
		video_pll_0_ref_clk_clk         : in    std_logic                     := '0';             --     video_pll_0_ref_clk.clk
		video_pll_0_ref_reset_reset     : in    std_logic                     := '0'              --   video_pll_0_ref_reset.reset
	);
end entity Computer_System;

architecture rtl of Computer_System is
	component Computer_System_ADC is
		generic (
			board          : string  := "DE10-Standard";
			board_rev      : string  := "Autodetect";
			tsclk          : integer := 0;
			numch          : integer := 0;
			max10pllmultby : integer := 0;
			max10plldivby  : integer := 0
		);
		port (
			clock       : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			address     : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			waitrequest : out std_logic;                                        -- waitrequest
			read        : in  std_logic                     := 'X';             -- read
			adc_sclk    : out std_logic;                                        -- export
			adc_cs_n    : out std_logic;                                        -- export
			adc_dout    : in  std_logic                     := 'X';             -- export
			adc_din     : out std_logic                                         -- export
		);
	end component Computer_System_ADC;

	component Computer_System_Arduino_GPIO is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			irq        : out   std_logic                                         -- irq
		);
	end component Computer_System_Arduino_GPIO;

	component Computer_System_Arduino_Reset_N is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component Computer_System_Arduino_Reset_N;

	component Computer_System_Expansion_JP1 is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic_vector(31 downto 0) := (others => 'X'); -- export
			irq        : out   std_logic                                         -- irq
		);
	end component Computer_System_Expansion_JP1;

	component Computer_System_HEX3_HEX0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component Computer_System_HEX3_HEX0;

	component Computer_System_Interval_Timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component Computer_System_Interval_Timer;

	component Computer_System_JTAG_UART is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component Computer_System_JTAG_UART;

	component Computer_System_JTAG_to_FPGA_Bridge is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component Computer_System_JTAG_to_FPGA_Bridge;

	component Computer_System_LEDs is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component Computer_System_LEDs;

	component Computer_System_Nios2 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			d_address                           : out std_logic_vector(31 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			E_ci_multi_done                     : in  std_logic                     := 'X';             -- done
			E_ci_multi_clk_en                   : out std_logic;                                        -- clk_en
			E_ci_multi_start                    : out std_logic;                                        -- start
			E_ci_result                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			D_ci_a                              : out std_logic_vector(4 downto 0);                     -- a
			D_ci_b                              : out std_logic_vector(4 downto 0);                     -- b
			D_ci_c                              : out std_logic_vector(4 downto 0);                     -- c
			D_ci_n                              : out std_logic_vector(7 downto 0);                     -- n
			D_ci_readra                         : out std_logic;                                        -- readra
			D_ci_readrb                         : out std_logic;                                        -- readrb
			D_ci_writerc                        : out std_logic;                                        -- writerc
			E_ci_dataa                          : out std_logic_vector(31 downto 0);                    -- dataa
			E_ci_datab                          : out std_logic_vector(31 downto 0);                    -- datab
			E_ci_multi_clock                    : out std_logic;                                        -- clk
			E_ci_multi_reset                    : out std_logic;                                        -- reset
			E_ci_multi_reset_req                : out std_logic;                                        -- reset_req
			W_ci_estatus                        : out std_logic;                                        -- estatus
			W_ci_ipending                       : out std_logic_vector(31 downto 0)                     -- ipending
		);
	end component Computer_System_Nios2;

	component fpoint_wrapper is
		generic (
			useDivider : integer := 0
		);
		port (
			clk    : in  std_logic                     := 'X';             -- clk
			clk_en : in  std_logic                     := 'X';             -- clk_en
			dataa  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			datab  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			n      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- n
			reset  : in  std_logic                     := 'X';             -- reset
			start  : in  std_logic                     := 'X';             -- start
			done   : out std_logic;                                        -- done
			result : out std_logic_vector(31 downto 0)                     -- result
		);
	end component fpoint_wrapper;

	component Computer_System_Onchip_SRAM is
		port (
			address     : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			address2    : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component Computer_System_Onchip_SRAM;

	component Computer_System_Pushbuttons is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component Computer_System_Pushbuttons;

	component Computer_System_SDRAM is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component Computer_System_SDRAM;

	component servo_control_port is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			rst        : in  std_logic                     := 'X';             -- reset
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			address    : in  std_logic                     := 'X';             -- address
			byteenable : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			control    : out std_logic                                         -- export
		);
	end component servo_control_port;

	component Computer_System_Slider_Switches is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(9 downto 0)  := (others => 'X')  -- export
		);
	end component Computer_System_Slider_Switches;

	component Computer_System_SysID is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component Computer_System_SysID;

	component Computer_System_System_PLL is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component Computer_System_System_PLL;

	component blinky_test_port is
		port (
			clk       : in  std_logic                    := 'X';             -- clk
			address   : in  std_logic                    := 'X';             -- address
			bytenable : in  std_logic                    := 'X';             -- byteenable
			write     : in  std_logic                    := 'X';             -- write
			read      : in  std_logic                    := 'X';             -- read
			writedata : in  std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			readdata  : out std_logic_vector(7 downto 0);                    -- readdata
			rst       : in  std_logic                    := 'X';             -- reset
			blinky    : out std_logic                                        -- export
		);
	end component blinky_test_port;

	component Computer_System_iServo0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(15 downto 0)                     -- export
		);
	end component Computer_System_iServo0;

	component Computer_System_video_lt24_controller_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			ready         : out std_logic;                                        -- ready
			startofpacket : in  std_logic                     := 'X';             -- startofpacket
			endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			data_in       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			data_in_valid : in  std_logic                     := 'X';             -- valid
			lt24_lcd_on   : out std_logic;                                        -- lcd_on
			lt24_reset_n  : out std_logic;                                        -- reset_n
			csx           : out std_logic;                                        -- csx
			data_to_lcd   : out std_logic_vector(15 downto 0);                    -- data
			rdx           : out std_logic;                                        -- rdx
			wrx           : out std_logic;                                        -- wrx
			data_not_cmd  : out std_logic                                         -- dcx
		);
	end component Computer_System_video_lt24_controller_0;

	component Computer_System_video_pixel_buffer_dma_0 is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic;                                        -- valid
			stream_data          : out std_logic_vector(15 downto 0)                     -- data
		);
	end component Computer_System_video_pixel_buffer_dma_0;

	component Computer_System_video_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			lcd_clk_clk        : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component Computer_System_video_pll_0;

	component altera_customins_master_translator is
		generic (
			SHARED_COMB_AND_MULTI : integer := 0
		);
		port (
			ci_slave_dataa            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result           : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n                : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra           : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb           : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc          : in  std_logic                     := 'X';             -- writerc
			ci_slave_a                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus          : in  std_logic                     := 'X';             -- estatus
			ci_slave_multi_clk        : in  std_logic                     := 'X';             -- clk
			ci_slave_multi_reset      : in  std_logic                     := 'X';             -- reset
			ci_slave_multi_clken      : in  std_logic                     := 'X';             -- clk_en
			ci_slave_multi_reset_req  : in  std_logic                     := 'X';             -- reset_req
			ci_slave_multi_start      : in  std_logic                     := 'X';             -- start
			ci_slave_multi_done       : out std_logic;                                        -- done
			comb_ci_master_dataa      : out std_logic_vector(31 downto 0);                    -- dataa
			comb_ci_master_datab      : out std_logic_vector(31 downto 0);                    -- datab
			comb_ci_master_result     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			comb_ci_master_n          : out std_logic_vector(7 downto 0);                     -- n
			comb_ci_master_readra     : out std_logic;                                        -- readra
			comb_ci_master_readrb     : out std_logic;                                        -- readrb
			comb_ci_master_writerc    : out std_logic;                                        -- writerc
			comb_ci_master_a          : out std_logic_vector(4 downto 0);                     -- a
			comb_ci_master_b          : out std_logic_vector(4 downto 0);                     -- b
			comb_ci_master_c          : out std_logic_vector(4 downto 0);                     -- c
			comb_ci_master_ipending   : out std_logic_vector(31 downto 0);                    -- ipending
			comb_ci_master_estatus    : out std_logic;                                        -- estatus
			multi_ci_master_clk       : out std_logic;                                        -- clk
			multi_ci_master_reset     : out std_logic;                                        -- reset
			multi_ci_master_clken     : out std_logic;                                        -- clk_en
			multi_ci_master_reset_req : out std_logic;                                        -- reset_req
			multi_ci_master_start     : out std_logic;                                        -- start
			multi_ci_master_done      : in  std_logic                     := 'X';             -- done
			multi_ci_master_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			multi_ci_master_datab     : out std_logic_vector(31 downto 0);                    -- datab
			multi_ci_master_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			multi_ci_master_n         : out std_logic_vector(7 downto 0);                     -- n
			multi_ci_master_readra    : out std_logic;                                        -- readra
			multi_ci_master_readrb    : out std_logic;                                        -- readrb
			multi_ci_master_writerc   : out std_logic;                                        -- writerc
			multi_ci_master_a         : out std_logic_vector(4 downto 0);                     -- a
			multi_ci_master_b         : out std_logic_vector(4 downto 0);                     -- b
			multi_ci_master_c         : out std_logic_vector(4 downto 0);                     -- c
			ci_slave_multi_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_dataa
			ci_slave_multi_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_datab
			ci_slave_multi_result     : out std_logic_vector(31 downto 0);                    -- multi_result
			ci_slave_multi_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- multi_n
			ci_slave_multi_readra     : in  std_logic                     := 'X';             -- multi_readra
			ci_slave_multi_readrb     : in  std_logic                     := 'X';             -- multi_readrb
			ci_slave_multi_writerc    : in  std_logic                     := 'X';             -- multi_writerc
			ci_slave_multi_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_a
			ci_slave_multi_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_b
			ci_slave_multi_c          : in  std_logic_vector(4 downto 0)  := (others => 'X')  -- multi_c
		);
	end component altera_customins_master_translator;

	component Computer_System_Nios2_custom_instruction_master_multi_xconnect is
		port (
			ci_slave_dataa       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result      : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra      : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb      : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc     : in  std_logic                     := 'X';             -- writerc
			ci_slave_a           : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b           : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c           : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus     : in  std_logic                     := 'X';             -- estatus
			ci_slave_clk         : in  std_logic                     := 'X';             -- clk
			ci_slave_reset       : in  std_logic                     := 'X';             -- reset
			ci_slave_clken       : in  std_logic                     := 'X';             -- clk_en
			ci_slave_reset_req   : in  std_logic                     := 'X';             -- reset_req
			ci_slave_start       : in  std_logic                     := 'X';             -- start
			ci_slave_done        : out std_logic;                                        -- done
			ci_master0_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master0_datab     : out std_logic_vector(31 downto 0);                    -- datab
			ci_master0_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master0_n         : out std_logic_vector(7 downto 0);                     -- n
			ci_master0_readra    : out std_logic;                                        -- readra
			ci_master0_readrb    : out std_logic;                                        -- readrb
			ci_master0_writerc   : out std_logic;                                        -- writerc
			ci_master0_a         : out std_logic_vector(4 downto 0);                     -- a
			ci_master0_b         : out std_logic_vector(4 downto 0);                     -- b
			ci_master0_c         : out std_logic_vector(4 downto 0);                     -- c
			ci_master0_ipending  : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master0_estatus   : out std_logic;                                        -- estatus
			ci_master0_clk       : out std_logic;                                        -- clk
			ci_master0_reset     : out std_logic;                                        -- reset
			ci_master0_clken     : out std_logic;                                        -- clk_en
			ci_master0_reset_req : out std_logic;                                        -- reset_req
			ci_master0_start     : out std_logic;                                        -- start
			ci_master0_done      : in  std_logic                     := 'X'              -- done
		);
	end component Computer_System_Nios2_custom_instruction_master_multi_xconnect;

	component altera_customins_slave_translator is
		generic (
			N_WIDTH          : integer := 8;
			USE_DONE         : integer := 1;
			NUM_FIXED_CYCLES : integer := 2
		);
		port (
			ci_slave_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result     : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra     : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb     : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc    : in  std_logic                     := 'X';             -- writerc
			ci_slave_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus    : in  std_logic                     := 'X';             -- estatus
			ci_slave_clk        : in  std_logic                     := 'X';             -- clk
			ci_slave_clken      : in  std_logic                     := 'X';             -- clk_en
			ci_slave_reset_req  : in  std_logic                     := 'X';             -- reset_req
			ci_slave_reset      : in  std_logic                     := 'X';             -- reset
			ci_slave_start      : in  std_logic                     := 'X';             -- start
			ci_slave_done       : out std_logic;                                        -- done
			ci_master_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master_datab     : out std_logic_vector(31 downto 0);                    -- datab
			ci_master_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master_n         : out std_logic_vector(1 downto 0);                     -- n
			ci_master_clk       : out std_logic;                                        -- clk
			ci_master_clken     : out std_logic;                                        -- clk_en
			ci_master_reset     : out std_logic;                                        -- reset
			ci_master_start     : out std_logic;                                        -- start
			ci_master_done      : in  std_logic                     := 'X';             -- done
			ci_master_readra    : out std_logic;                                        -- readra
			ci_master_readrb    : out std_logic;                                        -- readrb
			ci_master_writerc   : out std_logic;                                        -- writerc
			ci_master_a         : out std_logic_vector(4 downto 0);                     -- a
			ci_master_b         : out std_logic_vector(4 downto 0);                     -- b
			ci_master_c         : out std_logic_vector(4 downto 0);                     -- c
			ci_master_ipending  : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master_estatus   : out std_logic;                                        -- estatus
			ci_master_reset_req : out std_logic                                         -- reset_req
		);
	end component altera_customins_slave_translator;

	component Computer_System_mm_interconnect_0 is
		port (
			System_PLL_sys_clk_clk                                     : in  std_logic                     := 'X';             -- clk
			video_pll_0_lcd_clk_clk                                    : in  std_logic                     := 'X';             -- clk
			ADC_reset_reset_bridge_in_reset_reset                      : in  std_logic                     := 'X';             -- reset
			JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			Nios2_reset_reset_bridge_in_reset_reset                    : in  std_logic                     := 'X';             -- reset
			video_pixel_buffer_dma_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			JTAG_to_FPGA_Bridge_master_address                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			JTAG_to_FPGA_Bridge_master_waitrequest                     : out std_logic;                                        -- waitrequest
			JTAG_to_FPGA_Bridge_master_byteenable                      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			JTAG_to_FPGA_Bridge_master_read                            : in  std_logic                     := 'X';             -- read
			JTAG_to_FPGA_Bridge_master_readdata                        : out std_logic_vector(31 downto 0);                    -- readdata
			JTAG_to_FPGA_Bridge_master_readdatavalid                   : out std_logic;                                        -- readdatavalid
			JTAG_to_FPGA_Bridge_master_write                           : in  std_logic                     := 'X';             -- write
			JTAG_to_FPGA_Bridge_master_writedata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			Nios2_data_master_address                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			Nios2_data_master_waitrequest                              : out std_logic;                                        -- waitrequest
			Nios2_data_master_byteenable                               : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			Nios2_data_master_read                                     : in  std_logic                     := 'X';             -- read
			Nios2_data_master_readdata                                 : out std_logic_vector(31 downto 0);                    -- readdata
			Nios2_data_master_write                                    : in  std_logic                     := 'X';             -- write
			Nios2_data_master_writedata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			Nios2_data_master_debugaccess                              : in  std_logic                     := 'X';             -- debugaccess
			Nios2_instruction_master_address                           : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			Nios2_instruction_master_waitrequest                       : out std_logic;                                        -- waitrequest
			Nios2_instruction_master_read                              : in  std_logic                     := 'X';             -- read
			Nios2_instruction_master_readdata                          : out std_logic_vector(31 downto 0);                    -- readdata
			ADC_adc_slave_address                                      : out std_logic_vector(2 downto 0);                     -- address
			ADC_adc_slave_write                                        : out std_logic;                                        -- write
			ADC_adc_slave_read                                         : out std_logic;                                        -- read
			ADC_adc_slave_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ADC_adc_slave_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			ADC_adc_slave_waitrequest                                  : in  std_logic                     := 'X';             -- waitrequest
			Arduino_GPIO_s1_address                                    : out std_logic_vector(1 downto 0);                     -- address
			Arduino_GPIO_s1_write                                      : out std_logic;                                        -- write
			Arduino_GPIO_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Arduino_GPIO_s1_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			Arduino_GPIO_s1_chipselect                                 : out std_logic;                                        -- chipselect
			Arduino_Reset_N_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			Arduino_Reset_N_s1_write                                   : out std_logic;                                        -- write
			Arduino_Reset_N_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Arduino_Reset_N_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			Arduino_Reset_N_s1_chipselect                              : out std_logic;                                        -- chipselect
			blinky_test_0_avalon_slave_0_address                       : out std_logic_vector(0 downto 0);                     -- address
			blinky_test_0_avalon_slave_0_write                         : out std_logic;                                        -- write
			blinky_test_0_avalon_slave_0_read                          : out std_logic;                                        -- read
			blinky_test_0_avalon_slave_0_readdata                      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			blinky_test_0_avalon_slave_0_writedata                     : out std_logic_vector(7 downto 0);                     -- writedata
			blinky_test_0_avalon_slave_0_byteenable                    : out std_logic_vector(0 downto 0);                     -- byteenable
			Expansion_JP1_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			Expansion_JP1_s1_write                                     : out std_logic;                                        -- write
			Expansion_JP1_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Expansion_JP1_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			Expansion_JP1_s1_chipselect                                : out std_logic;                                        -- chipselect
			HEX3_HEX0_s1_address                                       : out std_logic_vector(1 downto 0);                     -- address
			HEX3_HEX0_s1_write                                         : out std_logic;                                        -- write
			HEX3_HEX0_s1_readdata                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX3_HEX0_s1_writedata                                     : out std_logic_vector(31 downto 0);                    -- writedata
			HEX3_HEX0_s1_chipselect                                    : out std_logic;                                        -- chipselect
			HEX5_HEX4_s1_address                                       : out std_logic_vector(1 downto 0);                     -- address
			HEX5_HEX4_s1_write                                         : out std_logic;                                        -- write
			HEX5_HEX4_s1_readdata                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX5_HEX4_s1_writedata                                     : out std_logic_vector(31 downto 0);                    -- writedata
			HEX5_HEX4_s1_chipselect                                    : out std_logic;                                        -- chipselect
			Interval_Timer_s1_address                                  : out std_logic_vector(2 downto 0);                     -- address
			Interval_Timer_s1_write                                    : out std_logic;                                        -- write
			Interval_Timer_s1_readdata                                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			Interval_Timer_s1_writedata                                : out std_logic_vector(15 downto 0);                    -- writedata
			Interval_Timer_s1_chipselect                               : out std_logic;                                        -- chipselect
			Interval_Timer_2_s1_address                                : out std_logic_vector(2 downto 0);                     -- address
			Interval_Timer_2_s1_write                                  : out std_logic;                                        -- write
			Interval_Timer_2_s1_readdata                               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			Interval_Timer_2_s1_writedata                              : out std_logic_vector(15 downto 0);                    -- writedata
			Interval_Timer_2_s1_chipselect                             : out std_logic;                                        -- chipselect
			iServo0_s1_address                                         : out std_logic_vector(1 downto 0);                     -- address
			iServo0_s1_write                                           : out std_logic;                                        -- write
			iServo0_s1_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			iServo0_s1_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			iServo0_s1_chipselect                                      : out std_logic;                                        -- chipselect
			iServo_0_s1_address                                        : out std_logic_vector(1 downto 0);                     -- address
			iServo_0_s1_write                                          : out std_logic;                                        -- write
			iServo_0_s1_readdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			iServo_0_s1_writedata                                      : out std_logic_vector(31 downto 0);                    -- writedata
			iServo_0_s1_chipselect                                     : out std_logic;                                        -- chipselect
			JTAG_UART_avalon_jtag_slave_address                        : out std_logic_vector(0 downto 0);                     -- address
			JTAG_UART_avalon_jtag_slave_write                          : out std_logic;                                        -- write
			JTAG_UART_avalon_jtag_slave_read                           : out std_logic;                                        -- read
			JTAG_UART_avalon_jtag_slave_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_UART_avalon_jtag_slave_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_UART_avalon_jtag_slave_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect                     : out std_logic;                                        -- chipselect
			LEDs_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			LEDs_s1_write                                              : out std_logic;                                        -- write
			LEDs_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LEDs_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			LEDs_s1_chipselect                                         : out std_logic;                                        -- chipselect
			Nios2_debug_mem_slave_address                              : out std_logic_vector(8 downto 0);                     -- address
			Nios2_debug_mem_slave_write                                : out std_logic;                                        -- write
			Nios2_debug_mem_slave_read                                 : out std_logic;                                        -- read
			Nios2_debug_mem_slave_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Nios2_debug_mem_slave_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			Nios2_debug_mem_slave_byteenable                           : out std_logic_vector(3 downto 0);                     -- byteenable
			Nios2_debug_mem_slave_waitrequest                          : in  std_logic                     := 'X';             -- waitrequest
			Nios2_debug_mem_slave_debugaccess                          : out std_logic;                                        -- debugaccess
			Onchip_SRAM_s1_address                                     : out std_logic_vector(13 downto 0);                    -- address
			Onchip_SRAM_s1_write                                       : out std_logic;                                        -- write
			Onchip_SRAM_s1_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Onchip_SRAM_s1_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			Onchip_SRAM_s1_byteenable                                  : out std_logic_vector(3 downto 0);                     -- byteenable
			Onchip_SRAM_s1_chipselect                                  : out std_logic;                                        -- chipselect
			Onchip_SRAM_s1_clken                                       : out std_logic;                                        -- clken
			Onchip_SRAM_s2_address                                     : out std_logic_vector(13 downto 0);                    -- address
			Onchip_SRAM_s2_write                                       : out std_logic;                                        -- write
			Onchip_SRAM_s2_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Onchip_SRAM_s2_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			Onchip_SRAM_s2_byteenable                                  : out std_logic_vector(3 downto 0);                     -- byteenable
			Onchip_SRAM_s2_chipselect                                  : out std_logic;                                        -- chipselect
			Onchip_SRAM_s2_clken                                       : out std_logic;                                        -- clken
			Pushbuttons_s1_address                                     : out std_logic_vector(1 downto 0);                     -- address
			Pushbuttons_s1_write                                       : out std_logic;                                        -- write
			Pushbuttons_s1_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Pushbuttons_s1_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			Pushbuttons_s1_chipselect                                  : out std_logic;                                        -- chipselect
			SDRAM_s1_address                                           : out std_logic_vector(24 downto 0);                    -- address
			SDRAM_s1_write                                             : out std_logic;                                        -- write
			SDRAM_s1_read                                              : out std_logic;                                        -- read
			SDRAM_s1_readdata                                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SDRAM_s1_writedata                                         : out std_logic_vector(15 downto 0);                    -- writedata
			SDRAM_s1_byteenable                                        : out std_logic_vector(1 downto 0);                     -- byteenable
			SDRAM_s1_readdatavalid                                     : in  std_logic                     := 'X';             -- readdatavalid
			SDRAM_s1_waitrequest                                       : in  std_logic                     := 'X';             -- waitrequest
			SDRAM_s1_chipselect                                        : out std_logic;                                        -- chipselect
			Servo0_servo_control_slave_address                         : out std_logic_vector(0 downto 0);                     -- address
			Servo0_servo_control_slave_write                           : out std_logic;                                        -- write
			Servo0_servo_control_slave_read                            : out std_logic;                                        -- read
			Servo0_servo_control_slave_readdata                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			Servo0_servo_control_slave_writedata                       : out std_logic_vector(15 downto 0);                    -- writedata
			Servo0_servo_control_slave_byteenable                      : out std_logic_vector(1 downto 0);                     -- byteenable
			Servo1_servo_control_slave_address                         : out std_logic_vector(0 downto 0);                     -- address
			Servo1_servo_control_slave_write                           : out std_logic;                                        -- write
			Servo1_servo_control_slave_read                            : out std_logic;                                        -- read
			Servo1_servo_control_slave_readdata                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			Servo1_servo_control_slave_writedata                       : out std_logic_vector(15 downto 0);                    -- writedata
			Servo1_servo_control_slave_byteenable                      : out std_logic_vector(1 downto 0);                     -- byteenable
			Slider_Switches_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			Slider_Switches_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SysID_control_slave_address                                : out std_logic_vector(0 downto 0);                     -- address
			SysID_control_slave_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			video_pixel_buffer_dma_0_avalon_control_slave_address      : out std_logic_vector(1 downto 0);                     -- address
			video_pixel_buffer_dma_0_avalon_control_slave_write        : out std_logic;                                        -- write
			video_pixel_buffer_dma_0_avalon_control_slave_read         : out std_logic;                                        -- read
			video_pixel_buffer_dma_0_avalon_control_slave_readdata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			video_pixel_buffer_dma_0_avalon_control_slave_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			video_pixel_buffer_dma_0_avalon_control_slave_byteenable   : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component Computer_System_mm_interconnect_0;

	component Computer_System_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Computer_System_irq_mapper;

	component computer_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component computer_system_rst_controller;

	component computer_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component computer_system_rst_controller_001;

	component computer_system_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component computer_system_rst_controller_002;

	signal video_pixel_buffer_dma_0_avalon_pixel_source_valid                         : std_logic;                     -- video_pixel_buffer_dma_0:stream_valid -> video_lt24_controller_0:data_in_valid
	signal video_pixel_buffer_dma_0_avalon_pixel_source_data                          : std_logic_vector(15 downto 0); -- video_pixel_buffer_dma_0:stream_data -> video_lt24_controller_0:data_in
	signal video_pixel_buffer_dma_0_avalon_pixel_source_ready                         : std_logic;                     -- video_lt24_controller_0:ready -> video_pixel_buffer_dma_0:stream_ready
	signal video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket                 : std_logic;                     -- video_pixel_buffer_dma_0:stream_startofpacket -> video_lt24_controller_0:startofpacket
	signal video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket                   : std_logic;                     -- video_pixel_buffer_dma_0:stream_endofpacket -> video_lt24_controller_0:endofpacket
	signal video_pll_0_lcd_clk_clk                                                    : std_logic;                     -- video_pll_0:lcd_clk_clk -> [mm_interconnect_0:video_pll_0_lcd_clk_clk, rst_controller_002:clk, video_lt24_controller_0:clk, video_pixel_buffer_dma_0:clk]
	signal system_pll_sys_clk_clk                                                     : std_logic;                     -- System_PLL:sys_clk_clk -> [ADC:clock, Arduino_GPIO:clk, Arduino_Reset_N:clk, Expansion_JP1:clk, HEX3_HEX0:clk, HEX5_HEX4:clk, Interval_Timer:clk, Interval_Timer_2:clk, JTAG_UART:clk, JTAG_UART_2nd_Core:clk, JTAG_to_FPGA_Bridge:clk_clk, LEDs:clk, Nios2:clk, Onchip_SRAM:clk, Pushbuttons:clk, SDRAM:clk, Servo0:clk, Servo1:clk, Slider_Switches:clk, SysID:clock, blinky_test_0:clk, iServo0:clk, iServo_0:clk, irq_mapper:clk, mm_interconnect_0:System_PLL_sys_clk_clk, rst_controller:clk, rst_controller_001:clk]
	signal system_pll_reset_source_reset                                              : std_logic;                     -- System_PLL:reset_source_reset -> [JTAG_to_FPGA_Bridge:clk_reset_reset, rst_controller:reset_in0, rst_controller_001:reset_in1]
	signal nios2_custom_instruction_master_readra                                     : std_logic;                     -- Nios2:D_ci_readra -> Nios2_custom_instruction_master_translator:ci_slave_readra
	signal nios2_custom_instruction_master_a                                          : std_logic_vector(4 downto 0);  -- Nios2:D_ci_a -> Nios2_custom_instruction_master_translator:ci_slave_a
	signal nios2_custom_instruction_master_b                                          : std_logic_vector(4 downto 0);  -- Nios2:D_ci_b -> Nios2_custom_instruction_master_translator:ci_slave_b
	signal nios2_custom_instruction_master_c                                          : std_logic_vector(4 downto 0);  -- Nios2:D_ci_c -> Nios2_custom_instruction_master_translator:ci_slave_c
	signal nios2_custom_instruction_master_readrb                                     : std_logic;                     -- Nios2:D_ci_readrb -> Nios2_custom_instruction_master_translator:ci_slave_readrb
	signal nios2_custom_instruction_master_clk                                        : std_logic;                     -- Nios2:E_ci_multi_clock -> Nios2_custom_instruction_master_translator:ci_slave_multi_clk
	signal nios2_custom_instruction_master_ipending                                   : std_logic_vector(31 downto 0); -- Nios2:W_ci_ipending -> Nios2_custom_instruction_master_translator:ci_slave_ipending
	signal nios2_custom_instruction_master_start                                      : std_logic;                     -- Nios2:E_ci_multi_start -> Nios2_custom_instruction_master_translator:ci_slave_multi_start
	signal nios2_custom_instruction_master_reset_req                                  : std_logic;                     -- Nios2:E_ci_multi_reset_req -> Nios2_custom_instruction_master_translator:ci_slave_multi_reset_req
	signal nios2_custom_instruction_master_done                                       : std_logic;                     -- Nios2_custom_instruction_master_translator:ci_slave_multi_done -> Nios2:E_ci_multi_done
	signal nios2_custom_instruction_master_n                                          : std_logic_vector(7 downto 0);  -- Nios2:D_ci_n -> Nios2_custom_instruction_master_translator:ci_slave_n
	signal nios2_custom_instruction_master_result                                     : std_logic_vector(31 downto 0); -- Nios2_custom_instruction_master_translator:ci_slave_result -> Nios2:E_ci_result
	signal nios2_custom_instruction_master_estatus                                    : std_logic;                     -- Nios2:W_ci_estatus -> Nios2_custom_instruction_master_translator:ci_slave_estatus
	signal nios2_custom_instruction_master_clk_en                                     : std_logic;                     -- Nios2:E_ci_multi_clk_en -> Nios2_custom_instruction_master_translator:ci_slave_multi_clken
	signal nios2_custom_instruction_master_datab                                      : std_logic_vector(31 downto 0); -- Nios2:E_ci_datab -> Nios2_custom_instruction_master_translator:ci_slave_datab
	signal nios2_custom_instruction_master_dataa                                      : std_logic_vector(31 downto 0); -- Nios2:E_ci_dataa -> Nios2_custom_instruction_master_translator:ci_slave_dataa
	signal nios2_custom_instruction_master_reset                                      : std_logic;                     -- Nios2:E_ci_multi_reset -> Nios2_custom_instruction_master_translator:ci_slave_multi_reset
	signal nios2_custom_instruction_master_writerc                                    : std_logic;                     -- Nios2:D_ci_writerc -> Nios2_custom_instruction_master_translator:ci_slave_writerc
	signal nios2_custom_instruction_master_translator_multi_ci_master_readra          : std_logic;                     -- Nios2_custom_instruction_master_translator:multi_ci_master_readra -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_readra
	signal nios2_custom_instruction_master_translator_multi_ci_master_a               : std_logic_vector(4 downto 0);  -- Nios2_custom_instruction_master_translator:multi_ci_master_a -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_a
	signal nios2_custom_instruction_master_translator_multi_ci_master_b               : std_logic_vector(4 downto 0);  -- Nios2_custom_instruction_master_translator:multi_ci_master_b -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_b
	signal nios2_custom_instruction_master_translator_multi_ci_master_clk             : std_logic;                     -- Nios2_custom_instruction_master_translator:multi_ci_master_clk -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_clk
	signal nios2_custom_instruction_master_translator_multi_ci_master_readrb          : std_logic;                     -- Nios2_custom_instruction_master_translator:multi_ci_master_readrb -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_readrb
	signal nios2_custom_instruction_master_translator_multi_ci_master_c               : std_logic_vector(4 downto 0);  -- Nios2_custom_instruction_master_translator:multi_ci_master_c -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_c
	signal nios2_custom_instruction_master_translator_multi_ci_master_start           : std_logic;                     -- Nios2_custom_instruction_master_translator:multi_ci_master_start -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_start
	signal nios2_custom_instruction_master_translator_multi_ci_master_reset_req       : std_logic;                     -- Nios2_custom_instruction_master_translator:multi_ci_master_reset_req -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	signal nios2_custom_instruction_master_translator_multi_ci_master_done            : std_logic;                     -- Nios2_custom_instruction_master_multi_xconnect:ci_slave_done -> Nios2_custom_instruction_master_translator:multi_ci_master_done
	signal nios2_custom_instruction_master_translator_multi_ci_master_n               : std_logic_vector(7 downto 0);  -- Nios2_custom_instruction_master_translator:multi_ci_master_n -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_n
	signal nios2_custom_instruction_master_translator_multi_ci_master_result          : std_logic_vector(31 downto 0); -- Nios2_custom_instruction_master_multi_xconnect:ci_slave_result -> Nios2_custom_instruction_master_translator:multi_ci_master_result
	signal nios2_custom_instruction_master_translator_multi_ci_master_clk_en          : std_logic;                     -- Nios2_custom_instruction_master_translator:multi_ci_master_clken -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_clken
	signal nios2_custom_instruction_master_translator_multi_ci_master_datab           : std_logic_vector(31 downto 0); -- Nios2_custom_instruction_master_translator:multi_ci_master_datab -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_datab
	signal nios2_custom_instruction_master_translator_multi_ci_master_dataa           : std_logic_vector(31 downto 0); -- Nios2_custom_instruction_master_translator:multi_ci_master_dataa -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_dataa
	signal nios2_custom_instruction_master_translator_multi_ci_master_reset           : std_logic;                     -- Nios2_custom_instruction_master_translator:multi_ci_master_reset -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_reset
	signal nios2_custom_instruction_master_translator_multi_ci_master_writerc         : std_logic;                     -- Nios2_custom_instruction_master_translator:multi_ci_master_writerc -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_writerc
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_readra           : std_logic;                     -- Nios2_custom_instruction_master_multi_xconnect:ci_master0_readra -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_a                : std_logic_vector(4 downto 0);  -- Nios2_custom_instruction_master_multi_xconnect:ci_master0_a -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_a
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_b                : std_logic_vector(4 downto 0);  -- Nios2_custom_instruction_master_multi_xconnect:ci_master0_b -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_b
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb           : std_logic;                     -- Nios2_custom_instruction_master_multi_xconnect:ci_master0_readrb -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_c                : std_logic_vector(4 downto 0);  -- Nios2_custom_instruction_master_multi_xconnect:ci_master0_c -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_c
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_clk              : std_logic;                     -- Nios2_custom_instruction_master_multi_xconnect:ci_master0_clk -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending         : std_logic_vector(31 downto 0); -- Nios2_custom_instruction_master_multi_xconnect:ci_master0_ipending -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_start            : std_logic;                     -- Nios2_custom_instruction_master_multi_xconnect:ci_master0_start -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_start
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req        : std_logic;                     -- Nios2_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_done             : std_logic;                     -- Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_done -> Nios2_custom_instruction_master_multi_xconnect:ci_master0_done
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_n                : std_logic_vector(7 downto 0);  -- Nios2_custom_instruction_master_multi_xconnect:ci_master0_n -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_n
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_result           : std_logic_vector(31 downto 0); -- Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_result -> Nios2_custom_instruction_master_multi_xconnect:ci_master0_result
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus          : std_logic;                     -- Nios2_custom_instruction_master_multi_xconnect:ci_master0_estatus -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en           : std_logic;                     -- Nios2_custom_instruction_master_multi_xconnect:ci_master0_clken -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_datab            : std_logic_vector(31 downto 0); -- Nios2_custom_instruction_master_multi_xconnect:ci_master0_datab -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa            : std_logic_vector(31 downto 0); -- Nios2_custom_instruction_master_multi_xconnect:ci_master0_dataa -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_reset            : std_logic;                     -- Nios2_custom_instruction_master_multi_xconnect:ci_master0_reset -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	signal nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc          : std_logic;                     -- Nios2_custom_instruction_master_multi_xconnect:ci_master0_writerc -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	signal nios2_custom_instruction_master_multi_slave_translator0_ci_master_result   : std_logic_vector(31 downto 0); -- Nios2_Floating_Point:result -> Nios2_custom_instruction_master_multi_slave_translator0:ci_master_result
	signal nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk      : std_logic;                     -- Nios2_custom_instruction_master_multi_slave_translator0:ci_master_clk -> Nios2_Floating_Point:clk
	signal nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en   : std_logic;                     -- Nios2_custom_instruction_master_multi_slave_translator0:ci_master_clken -> Nios2_Floating_Point:clk_en
	signal nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab    : std_logic_vector(31 downto 0); -- Nios2_custom_instruction_master_multi_slave_translator0:ci_master_datab -> Nios2_Floating_Point:datab
	signal nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa    : std_logic_vector(31 downto 0); -- Nios2_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> Nios2_Floating_Point:dataa
	signal nios2_custom_instruction_master_multi_slave_translator0_ci_master_start    : std_logic;                     -- Nios2_custom_instruction_master_multi_slave_translator0:ci_master_start -> Nios2_Floating_Point:start
	signal nios2_custom_instruction_master_multi_slave_translator0_ci_master_reset    : std_logic;                     -- Nios2_custom_instruction_master_multi_slave_translator0:ci_master_reset -> Nios2_Floating_Point:reset
	signal nios2_custom_instruction_master_multi_slave_translator0_ci_master_done     : std_logic;                     -- Nios2_Floating_Point:done -> Nios2_custom_instruction_master_multi_slave_translator0:ci_master_done
	signal nios2_custom_instruction_master_multi_slave_translator0_ci_master_n        : std_logic_vector(1 downto 0);  -- Nios2_custom_instruction_master_multi_slave_translator0:ci_master_n -> Nios2_Floating_Point:n
	signal nios2_data_master_readdata                                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:Nios2_data_master_readdata -> Nios2:d_readdata
	signal nios2_data_master_waitrequest                                              : std_logic;                     -- mm_interconnect_0:Nios2_data_master_waitrequest -> Nios2:d_waitrequest
	signal nios2_data_master_debugaccess                                              : std_logic;                     -- Nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Nios2_data_master_debugaccess
	signal nios2_data_master_address                                                  : std_logic_vector(31 downto 0); -- Nios2:d_address -> mm_interconnect_0:Nios2_data_master_address
	signal nios2_data_master_byteenable                                               : std_logic_vector(3 downto 0);  -- Nios2:d_byteenable -> mm_interconnect_0:Nios2_data_master_byteenable
	signal nios2_data_master_read                                                     : std_logic;                     -- Nios2:d_read -> mm_interconnect_0:Nios2_data_master_read
	signal nios2_data_master_write                                                    : std_logic;                     -- Nios2:d_write -> mm_interconnect_0:Nios2_data_master_write
	signal nios2_data_master_writedata                                                : std_logic_vector(31 downto 0); -- Nios2:d_writedata -> mm_interconnect_0:Nios2_data_master_writedata
	signal jtag_to_fpga_bridge_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_to_FPGA_Bridge_master_readdata -> JTAG_to_FPGA_Bridge:master_readdata
	signal jtag_to_fpga_bridge_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:JTAG_to_FPGA_Bridge_master_waitrequest -> JTAG_to_FPGA_Bridge:master_waitrequest
	signal jtag_to_fpga_bridge_master_address                                         : std_logic_vector(31 downto 0); -- JTAG_to_FPGA_Bridge:master_address -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_address
	signal jtag_to_fpga_bridge_master_read                                            : std_logic;                     -- JTAG_to_FPGA_Bridge:master_read -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_read
	signal jtag_to_fpga_bridge_master_byteenable                                      : std_logic_vector(3 downto 0);  -- JTAG_to_FPGA_Bridge:master_byteenable -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_byteenable
	signal jtag_to_fpga_bridge_master_readdatavalid                                   : std_logic;                     -- mm_interconnect_0:JTAG_to_FPGA_Bridge_master_readdatavalid -> JTAG_to_FPGA_Bridge:master_readdatavalid
	signal jtag_to_fpga_bridge_master_write                                           : std_logic;                     -- JTAG_to_FPGA_Bridge:master_write -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_write
	signal jtag_to_fpga_bridge_master_writedata                                       : std_logic_vector(31 downto 0); -- JTAG_to_FPGA_Bridge:master_writedata -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_writedata
	signal nios2_instruction_master_readdata                                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:Nios2_instruction_master_readdata -> Nios2:i_readdata
	signal nios2_instruction_master_waitrequest                                       : std_logic;                     -- mm_interconnect_0:Nios2_instruction_master_waitrequest -> Nios2:i_waitrequest
	signal nios2_instruction_master_address                                           : std_logic_vector(27 downto 0); -- Nios2:i_address -> mm_interconnect_0:Nios2_instruction_master_address
	signal nios2_instruction_master_read                                              : std_logic;                     -- Nios2:i_read -> mm_interconnect_0:Nios2_instruction_master_read
	signal mm_interconnect_0_adc_adc_slave_readdata                                   : std_logic_vector(31 downto 0); -- ADC:readdata -> mm_interconnect_0:ADC_adc_slave_readdata
	signal mm_interconnect_0_adc_adc_slave_waitrequest                                : std_logic;                     -- ADC:waitrequest -> mm_interconnect_0:ADC_adc_slave_waitrequest
	signal mm_interconnect_0_adc_adc_slave_address                                    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:ADC_adc_slave_address -> ADC:address
	signal mm_interconnect_0_adc_adc_slave_read                                       : std_logic;                     -- mm_interconnect_0:ADC_adc_slave_read -> ADC:read
	signal mm_interconnect_0_adc_adc_slave_write                                      : std_logic;                     -- mm_interconnect_0:ADC_adc_slave_write -> ADC:write
	signal mm_interconnect_0_adc_adc_slave_writedata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:ADC_adc_slave_writedata -> ADC:writedata
	signal mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata   : std_logic_vector(31 downto 0); -- video_pixel_buffer_dma_0:slave_readdata -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_readdata
	signal mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_address -> video_pixel_buffer_dma_0:slave_address
	signal mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read       : std_logic;                     -- mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_read -> video_pixel_buffer_dma_0:slave_read
	signal mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_byteenable -> video_pixel_buffer_dma_0:slave_byteenable
	signal mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write      : std_logic;                     -- mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_write -> video_pixel_buffer_dma_0:slave_write
	signal mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_writedata -> video_pixel_buffer_dma_0:slave_writedata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect                   : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata                     : std_logic_vector(31 downto 0); -- JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest                  : std_logic;                     -- JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address                      : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                         : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                        : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	signal mm_interconnect_0_blinky_test_0_avalon_slave_0_readdata                    : std_logic_vector(7 downto 0);  -- blinky_test_0:readdata -> mm_interconnect_0:blinky_test_0_avalon_slave_0_readdata
	signal mm_interconnect_0_blinky_test_0_avalon_slave_0_address                     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:blinky_test_0_avalon_slave_0_address -> blinky_test_0:address
	signal mm_interconnect_0_blinky_test_0_avalon_slave_0_read                        : std_logic;                     -- mm_interconnect_0:blinky_test_0_avalon_slave_0_read -> blinky_test_0:read
	signal mm_interconnect_0_blinky_test_0_avalon_slave_0_byteenable                  : std_logic_vector(0 downto 0);  -- mm_interconnect_0:blinky_test_0_avalon_slave_0_byteenable -> blinky_test_0:bytenable
	signal mm_interconnect_0_blinky_test_0_avalon_slave_0_write                       : std_logic;                     -- mm_interconnect_0:blinky_test_0_avalon_slave_0_write -> blinky_test_0:write
	signal mm_interconnect_0_blinky_test_0_avalon_slave_0_writedata                   : std_logic_vector(7 downto 0);  -- mm_interconnect_0:blinky_test_0_avalon_slave_0_writedata -> blinky_test_0:writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                             : std_logic_vector(31 downto 0); -- SysID:readdata -> mm_interconnect_0:SysID_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                              : std_logic_vector(0 downto 0);  -- mm_interconnect_0:SysID_control_slave_address -> SysID:address
	signal mm_interconnect_0_nios2_debug_mem_slave_readdata                           : std_logic_vector(31 downto 0); -- Nios2:debug_mem_slave_readdata -> mm_interconnect_0:Nios2_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_debug_mem_slave_waitrequest                        : std_logic;                     -- Nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:Nios2_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_debug_mem_slave_debugaccess                        : std_logic;                     -- mm_interconnect_0:Nios2_debug_mem_slave_debugaccess -> Nios2:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_debug_mem_slave_address                            : std_logic_vector(8 downto 0);  -- mm_interconnect_0:Nios2_debug_mem_slave_address -> Nios2:debug_mem_slave_address
	signal mm_interconnect_0_nios2_debug_mem_slave_read                               : std_logic;                     -- mm_interconnect_0:Nios2_debug_mem_slave_read -> Nios2:debug_mem_slave_read
	signal mm_interconnect_0_nios2_debug_mem_slave_byteenable                         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Nios2_debug_mem_slave_byteenable -> Nios2:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_debug_mem_slave_write                              : std_logic;                     -- mm_interconnect_0:Nios2_debug_mem_slave_write -> Nios2:debug_mem_slave_write
	signal mm_interconnect_0_nios2_debug_mem_slave_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:Nios2_debug_mem_slave_writedata -> Nios2:debug_mem_slave_writedata
	signal mm_interconnect_0_sdram_s1_chipselect                                      : std_logic;                     -- mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                                        : std_logic_vector(15 downto 0); -- SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                                     : std_logic;                     -- SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                                         : std_logic_vector(24 downto 0); -- mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	signal mm_interconnect_0_sdram_s1_read                                            : std_logic;                     -- mm_interconnect_0:SDRAM_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SDRAM_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                                   : std_logic;                     -- SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                                           : std_logic;                     -- mm_interconnect_0:SDRAM_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                                       : std_logic_vector(15 downto 0); -- mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	signal mm_interconnect_0_onchip_sram_s1_chipselect                                : std_logic;                     -- mm_interconnect_0:Onchip_SRAM_s1_chipselect -> Onchip_SRAM:chipselect
	signal mm_interconnect_0_onchip_sram_s1_readdata                                  : std_logic_vector(31 downto 0); -- Onchip_SRAM:readdata -> mm_interconnect_0:Onchip_SRAM_s1_readdata
	signal mm_interconnect_0_onchip_sram_s1_address                                   : std_logic_vector(13 downto 0); -- mm_interconnect_0:Onchip_SRAM_s1_address -> Onchip_SRAM:address
	signal mm_interconnect_0_onchip_sram_s1_byteenable                                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Onchip_SRAM_s1_byteenable -> Onchip_SRAM:byteenable
	signal mm_interconnect_0_onchip_sram_s1_write                                     : std_logic;                     -- mm_interconnect_0:Onchip_SRAM_s1_write -> Onchip_SRAM:write
	signal mm_interconnect_0_onchip_sram_s1_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:Onchip_SRAM_s1_writedata -> Onchip_SRAM:writedata
	signal mm_interconnect_0_onchip_sram_s1_clken                                     : std_logic;                     -- mm_interconnect_0:Onchip_SRAM_s1_clken -> Onchip_SRAM:clken
	signal mm_interconnect_0_leds_s1_chipselect                                       : std_logic;                     -- mm_interconnect_0:LEDs_s1_chipselect -> LEDs:chipselect
	signal mm_interconnect_0_leds_s1_readdata                                         : std_logic_vector(31 downto 0); -- LEDs:readdata -> mm_interconnect_0:LEDs_s1_readdata
	signal mm_interconnect_0_leds_s1_address                                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:LEDs_s1_address -> LEDs:address
	signal mm_interconnect_0_leds_s1_write                                            : std_logic;                     -- mm_interconnect_0:LEDs_s1_write -> mm_interconnect_0_leds_s1_write:in
	signal mm_interconnect_0_leds_s1_writedata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:LEDs_s1_writedata -> LEDs:writedata
	signal mm_interconnect_0_hex3_hex0_s1_chipselect                                  : std_logic;                     -- mm_interconnect_0:HEX3_HEX0_s1_chipselect -> HEX3_HEX0:chipselect
	signal mm_interconnect_0_hex3_hex0_s1_readdata                                    : std_logic_vector(31 downto 0); -- HEX3_HEX0:readdata -> mm_interconnect_0:HEX3_HEX0_s1_readdata
	signal mm_interconnect_0_hex3_hex0_s1_address                                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX3_HEX0_s1_address -> HEX3_HEX0:address
	signal mm_interconnect_0_hex3_hex0_s1_write                                       : std_logic;                     -- mm_interconnect_0:HEX3_HEX0_s1_write -> mm_interconnect_0_hex3_hex0_s1_write:in
	signal mm_interconnect_0_hex3_hex0_s1_writedata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX3_HEX0_s1_writedata -> HEX3_HEX0:writedata
	signal mm_interconnect_0_hex5_hex4_s1_chipselect                                  : std_logic;                     -- mm_interconnect_0:HEX5_HEX4_s1_chipselect -> HEX5_HEX4:chipselect
	signal mm_interconnect_0_hex5_hex4_s1_readdata                                    : std_logic_vector(31 downto 0); -- HEX5_HEX4:readdata -> mm_interconnect_0:HEX5_HEX4_s1_readdata
	signal mm_interconnect_0_hex5_hex4_s1_address                                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX5_HEX4_s1_address -> HEX5_HEX4:address
	signal mm_interconnect_0_hex5_hex4_s1_write                                       : std_logic;                     -- mm_interconnect_0:HEX5_HEX4_s1_write -> mm_interconnect_0_hex5_hex4_s1_write:in
	signal mm_interconnect_0_hex5_hex4_s1_writedata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX5_HEX4_s1_writedata -> HEX5_HEX4:writedata
	signal mm_interconnect_0_slider_switches_s1_readdata                              : std_logic_vector(31 downto 0); -- Slider_Switches:readdata -> mm_interconnect_0:Slider_Switches_s1_readdata
	signal mm_interconnect_0_slider_switches_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Slider_Switches_s1_address -> Slider_Switches:address
	signal mm_interconnect_0_pushbuttons_s1_chipselect                                : std_logic;                     -- mm_interconnect_0:Pushbuttons_s1_chipselect -> Pushbuttons:chipselect
	signal mm_interconnect_0_pushbuttons_s1_readdata                                  : std_logic_vector(31 downto 0); -- Pushbuttons:readdata -> mm_interconnect_0:Pushbuttons_s1_readdata
	signal mm_interconnect_0_pushbuttons_s1_address                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Pushbuttons_s1_address -> Pushbuttons:address
	signal mm_interconnect_0_pushbuttons_s1_write                                     : std_logic;                     -- mm_interconnect_0:Pushbuttons_s1_write -> mm_interconnect_0_pushbuttons_s1_write:in
	signal mm_interconnect_0_pushbuttons_s1_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:Pushbuttons_s1_writedata -> Pushbuttons:writedata
	signal mm_interconnect_0_expansion_jp1_s1_chipselect                              : std_logic;                     -- mm_interconnect_0:Expansion_JP1_s1_chipselect -> Expansion_JP1:chipselect
	signal mm_interconnect_0_expansion_jp1_s1_readdata                                : std_logic_vector(31 downto 0); -- Expansion_JP1:readdata -> mm_interconnect_0:Expansion_JP1_s1_readdata
	signal mm_interconnect_0_expansion_jp1_s1_address                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Expansion_JP1_s1_address -> Expansion_JP1:address
	signal mm_interconnect_0_expansion_jp1_s1_write                                   : std_logic;                     -- mm_interconnect_0:Expansion_JP1_s1_write -> mm_interconnect_0_expansion_jp1_s1_write:in
	signal mm_interconnect_0_expansion_jp1_s1_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:Expansion_JP1_s1_writedata -> Expansion_JP1:writedata
	signal mm_interconnect_0_arduino_gpio_s1_chipselect                               : std_logic;                     -- mm_interconnect_0:Arduino_GPIO_s1_chipselect -> Arduino_GPIO:chipselect
	signal mm_interconnect_0_arduino_gpio_s1_readdata                                 : std_logic_vector(31 downto 0); -- Arduino_GPIO:readdata -> mm_interconnect_0:Arduino_GPIO_s1_readdata
	signal mm_interconnect_0_arduino_gpio_s1_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Arduino_GPIO_s1_address -> Arduino_GPIO:address
	signal mm_interconnect_0_arduino_gpio_s1_write                                    : std_logic;                     -- mm_interconnect_0:Arduino_GPIO_s1_write -> mm_interconnect_0_arduino_gpio_s1_write:in
	signal mm_interconnect_0_arduino_gpio_s1_writedata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:Arduino_GPIO_s1_writedata -> Arduino_GPIO:writedata
	signal mm_interconnect_0_arduino_reset_n_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:Arduino_Reset_N_s1_chipselect -> Arduino_Reset_N:chipselect
	signal mm_interconnect_0_arduino_reset_n_s1_readdata                              : std_logic_vector(31 downto 0); -- Arduino_Reset_N:readdata -> mm_interconnect_0:Arduino_Reset_N_s1_readdata
	signal mm_interconnect_0_arduino_reset_n_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Arduino_Reset_N_s1_address -> Arduino_Reset_N:address
	signal mm_interconnect_0_arduino_reset_n_s1_write                                 : std_logic;                     -- mm_interconnect_0:Arduino_Reset_N_s1_write -> mm_interconnect_0_arduino_reset_n_s1_write:in
	signal mm_interconnect_0_arduino_reset_n_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:Arduino_Reset_N_s1_writedata -> Arduino_Reset_N:writedata
	signal mm_interconnect_0_interval_timer_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:Interval_Timer_s1_chipselect -> Interval_Timer:chipselect
	signal mm_interconnect_0_interval_timer_s1_readdata                               : std_logic_vector(15 downto 0); -- Interval_Timer:readdata -> mm_interconnect_0:Interval_Timer_s1_readdata
	signal mm_interconnect_0_interval_timer_s1_address                                : std_logic_vector(2 downto 0);  -- mm_interconnect_0:Interval_Timer_s1_address -> Interval_Timer:address
	signal mm_interconnect_0_interval_timer_s1_write                                  : std_logic;                     -- mm_interconnect_0:Interval_Timer_s1_write -> mm_interconnect_0_interval_timer_s1_write:in
	signal mm_interconnect_0_interval_timer_s1_writedata                              : std_logic_vector(15 downto 0); -- mm_interconnect_0:Interval_Timer_s1_writedata -> Interval_Timer:writedata
	signal mm_interconnect_0_interval_timer_2_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:Interval_Timer_2_s1_chipselect -> Interval_Timer_2:chipselect
	signal mm_interconnect_0_interval_timer_2_s1_readdata                             : std_logic_vector(15 downto 0); -- Interval_Timer_2:readdata -> mm_interconnect_0:Interval_Timer_2_s1_readdata
	signal mm_interconnect_0_interval_timer_2_s1_address                              : std_logic_vector(2 downto 0);  -- mm_interconnect_0:Interval_Timer_2_s1_address -> Interval_Timer_2:address
	signal mm_interconnect_0_interval_timer_2_s1_write                                : std_logic;                     -- mm_interconnect_0:Interval_Timer_2_s1_write -> mm_interconnect_0_interval_timer_2_s1_write:in
	signal mm_interconnect_0_interval_timer_2_s1_writedata                            : std_logic_vector(15 downto 0); -- mm_interconnect_0:Interval_Timer_2_s1_writedata -> Interval_Timer_2:writedata
	signal mm_interconnect_0_iservo0_s1_chipselect                                    : std_logic;                     -- mm_interconnect_0:iServo0_s1_chipselect -> iServo0:chipselect
	signal mm_interconnect_0_iservo0_s1_readdata                                      : std_logic_vector(31 downto 0); -- iServo0:readdata -> mm_interconnect_0:iServo0_s1_readdata
	signal mm_interconnect_0_iservo0_s1_address                                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:iServo0_s1_address -> iServo0:address
	signal mm_interconnect_0_iservo0_s1_write                                         : std_logic;                     -- mm_interconnect_0:iServo0_s1_write -> mm_interconnect_0_iservo0_s1_write:in
	signal mm_interconnect_0_iservo0_s1_writedata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:iServo0_s1_writedata -> iServo0:writedata
	signal mm_interconnect_0_iservo_0_s1_chipselect                                   : std_logic;                     -- mm_interconnect_0:iServo_0_s1_chipselect -> iServo_0:chipselect
	signal mm_interconnect_0_iservo_0_s1_readdata                                     : std_logic_vector(31 downto 0); -- iServo_0:readdata -> mm_interconnect_0:iServo_0_s1_readdata
	signal mm_interconnect_0_iservo_0_s1_address                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:iServo_0_s1_address -> iServo_0:address
	signal mm_interconnect_0_iservo_0_s1_write                                        : std_logic;                     -- mm_interconnect_0:iServo_0_s1_write -> mm_interconnect_0_iservo_0_s1_write:in
	signal mm_interconnect_0_iservo_0_s1_writedata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:iServo_0_s1_writedata -> iServo_0:writedata
	signal mm_interconnect_0_servo0_servo_control_slave_readdata                      : std_logic_vector(15 downto 0); -- Servo0:readdata -> mm_interconnect_0:Servo0_servo_control_slave_readdata
	signal mm_interconnect_0_servo0_servo_control_slave_address                       : std_logic_vector(0 downto 0);  -- mm_interconnect_0:Servo0_servo_control_slave_address -> Servo0:address
	signal mm_interconnect_0_servo0_servo_control_slave_read                          : std_logic;                     -- mm_interconnect_0:Servo0_servo_control_slave_read -> Servo0:read
	signal mm_interconnect_0_servo0_servo_control_slave_byteenable                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Servo0_servo_control_slave_byteenable -> Servo0:byteenable
	signal mm_interconnect_0_servo0_servo_control_slave_write                         : std_logic;                     -- mm_interconnect_0:Servo0_servo_control_slave_write -> Servo0:write
	signal mm_interconnect_0_servo0_servo_control_slave_writedata                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:Servo0_servo_control_slave_writedata -> Servo0:writedata
	signal mm_interconnect_0_servo1_servo_control_slave_readdata                      : std_logic_vector(15 downto 0); -- Servo1:readdata -> mm_interconnect_0:Servo1_servo_control_slave_readdata
	signal mm_interconnect_0_servo1_servo_control_slave_address                       : std_logic_vector(0 downto 0);  -- mm_interconnect_0:Servo1_servo_control_slave_address -> Servo1:address
	signal mm_interconnect_0_servo1_servo_control_slave_read                          : std_logic;                     -- mm_interconnect_0:Servo1_servo_control_slave_read -> Servo1:read
	signal mm_interconnect_0_servo1_servo_control_slave_byteenable                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Servo1_servo_control_slave_byteenable -> Servo1:byteenable
	signal mm_interconnect_0_servo1_servo_control_slave_write                         : std_logic;                     -- mm_interconnect_0:Servo1_servo_control_slave_write -> Servo1:write
	signal mm_interconnect_0_servo1_servo_control_slave_writedata                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:Servo1_servo_control_slave_writedata -> Servo1:writedata
	signal mm_interconnect_0_onchip_sram_s2_chipselect                                : std_logic;                     -- mm_interconnect_0:Onchip_SRAM_s2_chipselect -> Onchip_SRAM:chipselect2
	signal mm_interconnect_0_onchip_sram_s2_readdata                                  : std_logic_vector(31 downto 0); -- Onchip_SRAM:readdata2 -> mm_interconnect_0:Onchip_SRAM_s2_readdata
	signal mm_interconnect_0_onchip_sram_s2_address                                   : std_logic_vector(13 downto 0); -- mm_interconnect_0:Onchip_SRAM_s2_address -> Onchip_SRAM:address2
	signal mm_interconnect_0_onchip_sram_s2_byteenable                                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Onchip_SRAM_s2_byteenable -> Onchip_SRAM:byteenable2
	signal mm_interconnect_0_onchip_sram_s2_write                                     : std_logic;                     -- mm_interconnect_0:Onchip_SRAM_s2_write -> Onchip_SRAM:write2
	signal mm_interconnect_0_onchip_sram_s2_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:Onchip_SRAM_s2_writedata -> Onchip_SRAM:writedata2
	signal mm_interconnect_0_onchip_sram_s2_clken                                     : std_logic;                     -- mm_interconnect_0:Onchip_SRAM_s2_clken -> Onchip_SRAM:clken2
	signal irq_mapper_receiver0_irq                                                   : std_logic;                     -- Pushbuttons:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                   : std_logic;                     -- Expansion_JP1:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                   : std_logic;                     -- Arduino_GPIO:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                                   : std_logic;                     -- JTAG_UART:av_irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                                   : std_logic;                     -- Interval_Timer:irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                                   : std_logic;                     -- Interval_Timer_2:irq -> irq_mapper:receiver5_irq
	signal nios2_irq_irq                                                              : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> Nios2:irq
	signal rst_controller_reset_out_reset                                             : std_logic;                     -- rst_controller:reset_out -> [ADC:reset, Onchip_SRAM:reset, Servo0:rst, Servo1:rst, blinky_test_0:rst, mm_interconnect_0:ADC_reset_reset_bridge_in_reset_reset, mm_interconnect_0:JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                         : std_logic;                     -- rst_controller:reset_req -> [Onchip_SRAM:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                                         : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:Nios2_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal nios2_debug_reset_request_reset                                            : std_logic;                     -- Nios2:debug_reset_request -> rst_controller_001:reset_in0
	signal rst_controller_002_reset_out_reset                                         : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:video_pixel_buffer_dma_0_reset_reset_bridge_in_reset_reset, video_lt24_controller_0:reset, video_pixel_buffer_dma_0:reset]
	signal video_pll_0_reset_source_reset                                             : std_logic;                     -- video_pll_0:reset_source_reset -> rst_controller_002:reset_in0
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv               : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> JTAG_UART:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv              : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> JTAG_UART:av_write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                                  : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> SDRAM:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> SDRAM:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                                 : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> SDRAM:az_wr_n
	signal mm_interconnect_0_leds_s1_write_ports_inv                                  : std_logic;                     -- mm_interconnect_0_leds_s1_write:inv -> LEDs:write_n
	signal mm_interconnect_0_hex3_hex0_s1_write_ports_inv                             : std_logic;                     -- mm_interconnect_0_hex3_hex0_s1_write:inv -> HEX3_HEX0:write_n
	signal mm_interconnect_0_hex5_hex4_s1_write_ports_inv                             : std_logic;                     -- mm_interconnect_0_hex5_hex4_s1_write:inv -> HEX5_HEX4:write_n
	signal mm_interconnect_0_pushbuttons_s1_write_ports_inv                           : std_logic;                     -- mm_interconnect_0_pushbuttons_s1_write:inv -> Pushbuttons:write_n
	signal mm_interconnect_0_expansion_jp1_s1_write_ports_inv                         : std_logic;                     -- mm_interconnect_0_expansion_jp1_s1_write:inv -> Expansion_JP1:write_n
	signal mm_interconnect_0_arduino_gpio_s1_write_ports_inv                          : std_logic;                     -- mm_interconnect_0_arduino_gpio_s1_write:inv -> Arduino_GPIO:write_n
	signal mm_interconnect_0_arduino_reset_n_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_0_arduino_reset_n_s1_write:inv -> Arduino_Reset_N:write_n
	signal mm_interconnect_0_interval_timer_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_interval_timer_s1_write:inv -> Interval_Timer:write_n
	signal mm_interconnect_0_interval_timer_2_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_interval_timer_2_s1_write:inv -> Interval_Timer_2:write_n
	signal mm_interconnect_0_iservo0_s1_write_ports_inv                               : std_logic;                     -- mm_interconnect_0_iservo0_s1_write:inv -> iServo0:write_n
	signal mm_interconnect_0_iservo_0_s1_write_ports_inv                              : std_logic;                     -- mm_interconnect_0_iservo_0_s1_write:inv -> iServo_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                                   : std_logic;                     -- rst_controller_reset_out_reset:inv -> [Arduino_GPIO:reset_n, Arduino_Reset_N:reset_n, Expansion_JP1:reset_n, HEX3_HEX0:reset_n, HEX5_HEX4:reset_n, Interval_Timer:reset_n, Interval_Timer_2:reset_n, JTAG_UART:rst_n, JTAG_UART_2nd_Core:rst_n, LEDs:reset_n, Pushbuttons:reset_n, SDRAM:reset_n, Slider_Switches:reset_n, SysID:reset_n, iServo0:reset_n, iServo_0:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                               : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> Nios2:reset_n

begin

	adc : component Computer_System_ADC
		generic map (
			board          => "DE10-Lite",
			board_rev      => "Autodetect",
			tsclk          => 10,
			numch          => 5,
			max10pllmultby => 1,
			max10plldivby  => 10
		)
		port map (
			clock       => system_pll_sys_clk_clk,                      --       clk.clk
			reset       => rst_controller_reset_out_reset,              --     reset.reset
			write       => mm_interconnect_0_adc_adc_slave_write,       -- adc_slave.write
			readdata    => mm_interconnect_0_adc_adc_slave_readdata,    --          .readdata
			writedata   => mm_interconnect_0_adc_adc_slave_writedata,   --          .writedata
			address     => mm_interconnect_0_adc_adc_slave_address,     --          .address
			waitrequest => mm_interconnect_0_adc_adc_slave_waitrequest, --          .waitrequest
			read        => mm_interconnect_0_adc_adc_slave_read,        --          .read
			adc_sclk    => open,                                        -- (terminated)
			adc_cs_n    => open,                                        -- (terminated)
			adc_dout    => '0',                                         -- (terminated)
			adc_din     => open                                         -- (terminated)
		);

	arduino_gpio : component Computer_System_Arduino_GPIO
		port map (
			clk        => system_pll_sys_clk_clk,                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_0_arduino_gpio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_arduino_gpio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_arduino_gpio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_arduino_gpio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_arduino_gpio_s1_readdata,        --                    .readdata
			bidir_port => arduino_gpio_export,                               -- external_connection.export
			irq        => irq_mapper_receiver2_irq                           --                 irq.irq
		);

	arduino_reset_n : component Computer_System_Arduino_Reset_N
		port map (
			clk        => system_pll_sys_clk_clk,                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,             --               reset.reset_n
			address    => mm_interconnect_0_arduino_reset_n_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_arduino_reset_n_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_arduino_reset_n_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_arduino_reset_n_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_arduino_reset_n_s1_readdata,        --                    .readdata
			out_port   => arduino_reset_n_export                                -- external_connection.export
		);

	expansion_jp1 : component Computer_System_Expansion_JP1
		port map (
			clk        => system_pll_sys_clk_clk,                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           --               reset.reset_n
			address    => mm_interconnect_0_expansion_jp1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_expansion_jp1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_expansion_jp1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_expansion_jp1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_expansion_jp1_s1_readdata,        --                    .readdata
			bidir_port => expansion_jp1_export,                               -- external_connection.export
			irq        => irq_mapper_receiver1_irq                            --                 irq.irq
		);

	hex3_hex0 : component Computer_System_HEX3_HEX0
		port map (
			clk        => system_pll_sys_clk_clk,                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_hex3_hex0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex3_hex0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex3_hex0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex3_hex0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex3_hex0_s1_readdata,        --                    .readdata
			out_port   => hex3_hex0_export                                -- external_connection.export
		);

	hex5_hex4 : component Computer_System_HEX3_HEX0
		port map (
			clk        => system_pll_sys_clk_clk,                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_hex5_hex4_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex5_hex4_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex5_hex4_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex5_hex4_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex5_hex4_s1_readdata,        --                    .readdata
			out_port   => hex5_hex4_export                                -- external_connection.export
		);

	interval_timer : component Computer_System_Interval_Timer
		port map (
			clk        => system_pll_sys_clk_clk,                              --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,            -- reset.reset_n
			address    => mm_interconnect_0_interval_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_interval_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_interval_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_interval_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_interval_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver4_irq                             --   irq.irq
		);

	interval_timer_2 : component Computer_System_Interval_Timer
		port map (
			clk        => system_pll_sys_clk_clk,                                --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              -- reset.reset_n
			address    => mm_interconnect_0_interval_timer_2_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_interval_timer_2_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_interval_timer_2_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_interval_timer_2_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_interval_timer_2_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver5_irq                               --   irq.irq
		);

	jtag_uart : component Computer_System_JTAG_UART
		port map (
			clk            => system_pll_sys_clk_clk,                                        --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver3_irq                                       --               irq.irq
		);

	jtag_uart_2nd_core : component Computer_System_JTAG_UART
		port map (
			clk            => system_pll_sys_clk_clk,                   --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv, --             reset.reset_n
			av_chipselect  => open,                                     -- avalon_jtag_slave.chipselect
			av_address     => open,                                     --                  .address
			av_read_n      => open,                                     --                  .read_n
			av_readdata    => open,                                     --                  .readdata
			av_write_n     => open,                                     --                  .write_n
			av_writedata   => open,                                     --                  .writedata
			av_waitrequest => open,                                     --                  .waitrequest
			av_irq         => open                                      --               irq.irq
		);

	jtag_to_fpga_bridge : component Computer_System_JTAG_to_FPGA_Bridge
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => system_pll_sys_clk_clk,                   --          clk.clk
			clk_reset_reset      => system_pll_reset_source_reset,            --    clk_reset.reset
			master_address       => jtag_to_fpga_bridge_master_address,       --       master.address
			master_readdata      => jtag_to_fpga_bridge_master_readdata,      --             .readdata
			master_read          => jtag_to_fpga_bridge_master_read,          --             .read
			master_write         => jtag_to_fpga_bridge_master_write,         --             .write
			master_writedata     => jtag_to_fpga_bridge_master_writedata,     --             .writedata
			master_waitrequest   => jtag_to_fpga_bridge_master_waitrequest,   --             .waitrequest
			master_readdatavalid => jtag_to_fpga_bridge_master_readdatavalid, --             .readdatavalid
			master_byteenable    => jtag_to_fpga_bridge_master_byteenable,    --             .byteenable
			master_reset_reset   => open                                      -- master_reset.reset
		);

	leds : component Computer_System_LEDs
		port map (
			clk        => system_pll_sys_clk_clk,                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_leds_s1_readdata,        --                    .readdata
			out_port   => leds_export                                -- external_connection.export
		);

	nios2 : component Computer_System_Nios2
		port map (
			clk                                 => system_pll_sys_clk_clk,                              --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,        --                     reset.reset_n
			d_address                           => nios2_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_data_master_read,                              --                          .read
			d_readdata                          => nios2_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_data_master_write,                             --                          .write
			d_writedata                         => nios2_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_debug_mem_slave_writedata,   --                          .writedata
			E_ci_multi_done                     => nios2_custom_instruction_master_done,                -- custom_instruction_master.done
			E_ci_multi_clk_en                   => nios2_custom_instruction_master_clk_en,              --                          .clk_en
			E_ci_multi_start                    => nios2_custom_instruction_master_start,               --                          .start
			E_ci_result                         => nios2_custom_instruction_master_result,              --                          .result
			D_ci_a                              => nios2_custom_instruction_master_a,                   --                          .a
			D_ci_b                              => nios2_custom_instruction_master_b,                   --                          .b
			D_ci_c                              => nios2_custom_instruction_master_c,                   --                          .c
			D_ci_n                              => nios2_custom_instruction_master_n,                   --                          .n
			D_ci_readra                         => nios2_custom_instruction_master_readra,              --                          .readra
			D_ci_readrb                         => nios2_custom_instruction_master_readrb,              --                          .readrb
			D_ci_writerc                        => nios2_custom_instruction_master_writerc,             --                          .writerc
			E_ci_dataa                          => nios2_custom_instruction_master_dataa,               --                          .dataa
			E_ci_datab                          => nios2_custom_instruction_master_datab,               --                          .datab
			E_ci_multi_clock                    => nios2_custom_instruction_master_clk,                 --                          .clk
			E_ci_multi_reset                    => nios2_custom_instruction_master_reset,               --                          .reset
			E_ci_multi_reset_req                => nios2_custom_instruction_master_reset_req,           --                          .reset_req
			W_ci_estatus                        => nios2_custom_instruction_master_estatus,             --                          .estatus
			W_ci_ipending                       => nios2_custom_instruction_master_ipending             --                          .ipending
		);

	nios2_floating_point : component fpoint_wrapper
		generic map (
			useDivider => 1
		)
		port map (
			clk    => nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk,    -- s1.clk
			clk_en => nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en, --   .clk_en
			dataa  => nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa,  --   .dataa
			datab  => nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab,  --   .datab
			n      => nios2_custom_instruction_master_multi_slave_translator0_ci_master_n,      --   .n
			reset  => nios2_custom_instruction_master_multi_slave_translator0_ci_master_reset,  --   .reset
			start  => nios2_custom_instruction_master_multi_slave_translator0_ci_master_start,  --   .start
			done   => nios2_custom_instruction_master_multi_slave_translator0_ci_master_done,   --   .done
			result => nios2_custom_instruction_master_multi_slave_translator0_ci_master_result  --   .result
		);

	onchip_sram : component Computer_System_Onchip_SRAM
		port map (
			address     => mm_interconnect_0_onchip_sram_s1_address,    --     s1.address
			clken       => mm_interconnect_0_onchip_sram_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_onchip_sram_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_onchip_sram_s1_write,      --       .write
			readdata    => mm_interconnect_0_onchip_sram_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_onchip_sram_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_onchip_sram_s1_byteenable, --       .byteenable
			address2    => mm_interconnect_0_onchip_sram_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_0_onchip_sram_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_0_onchip_sram_s2_clken,      --       .clken
			write2      => mm_interconnect_0_onchip_sram_s2_write,      --       .write
			readdata2   => mm_interconnect_0_onchip_sram_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_0_onchip_sram_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_0_onchip_sram_s2_byteenable, --       .byteenable
			clk         => system_pll_sys_clk_clk,                      --   clk1.clk
			reset       => rst_controller_reset_out_reset,              -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,          --       .reset_req
			freeze      => '0'                                          -- (terminated)
		);

	pushbuttons : component Computer_System_Pushbuttons
		port map (
			clk        => system_pll_sys_clk_clk,                           --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_pushbuttons_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pushbuttons_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pushbuttons_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pushbuttons_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pushbuttons_s1_readdata,        --                    .readdata
			in_port    => pushbuttons_export,                               -- external_connection.export
			irq        => irq_mapper_receiver0_irq                          --                 irq.irq
		);

	sdram : component Computer_System_SDRAM
		port map (
			clk            => system_pll_sys_clk_clk,                          --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	servo0 : component servo_control_port
		port map (
			clk        => system_pll_sys_clk_clk,                                  --                 clk.clk
			rst        => rst_controller_reset_out_reset,                          --                 rst.reset
			readdata   => mm_interconnect_0_servo0_servo_control_slave_readdata,   -- servo_control_slave.readdata
			writedata  => mm_interconnect_0_servo0_servo_control_slave_writedata,  --                    .writedata
			read       => mm_interconnect_0_servo0_servo_control_slave_read,       --                    .read
			write      => mm_interconnect_0_servo0_servo_control_slave_write,      --                    .write
			address    => mm_interconnect_0_servo0_servo_control_slave_address(0), --                    .address
			byteenable => mm_interconnect_0_servo0_servo_control_slave_byteenable, --                    .byteenable
			control    => servo_control_0_export                                   -- external_connection.export
		);

	servo1 : component servo_control_port
		port map (
			clk        => system_pll_sys_clk_clk,                                  --                 clk.clk
			rst        => rst_controller_reset_out_reset,                          --                 rst.reset
			readdata   => mm_interconnect_0_servo1_servo_control_slave_readdata,   -- servo_control_slave.readdata
			writedata  => mm_interconnect_0_servo1_servo_control_slave_writedata,  --                    .writedata
			read       => mm_interconnect_0_servo1_servo_control_slave_read,       --                    .read
			write      => mm_interconnect_0_servo1_servo_control_slave_write,      --                    .write
			address    => mm_interconnect_0_servo1_servo_control_slave_address(0), --                    .address
			byteenable => mm_interconnect_0_servo1_servo_control_slave_byteenable, --                    .byteenable
			control    => servo_control_1_export                                   -- external_connection.export
		);

	slider_switches : component Computer_System_Slider_Switches
		port map (
			clk      => system_pll_sys_clk_clk,                        --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address  => mm_interconnect_0_slider_switches_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_slider_switches_s1_readdata, --                    .readdata
			in_port  => slider_switches_export                         -- external_connection.export
		);

	sysid : component Computer_System_SysID
		port map (
			clock    => system_pll_sys_clk_clk,                           --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	system_pll : component Computer_System_System_PLL
		port map (
			ref_clk_clk        => system_pll_ref_clk_clk,        --      ref_clk.clk
			ref_reset_reset    => system_pll_ref_reset_reset,    --    ref_reset.reset
			sys_clk_clk        => system_pll_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => sdram_clk_clk,                 --    sdram_clk.clk
			reset_source_reset => system_pll_reset_source_reset  -- reset_source.reset
		);

	blinky_test_0 : component blinky_test_port
		port map (
			clk       => system_pll_sys_clk_clk,                                       --          clock.clk
			address   => mm_interconnect_0_blinky_test_0_avalon_slave_0_address(0),    -- avalon_slave_0.address
			bytenable => mm_interconnect_0_blinky_test_0_avalon_slave_0_byteenable(0), --               .byteenable
			write     => mm_interconnect_0_blinky_test_0_avalon_slave_0_write,         --               .write
			read      => mm_interconnect_0_blinky_test_0_avalon_slave_0_read,          --               .read
			writedata => mm_interconnect_0_blinky_test_0_avalon_slave_0_writedata,     --               .writedata
			readdata  => mm_interconnect_0_blinky_test_0_avalon_slave_0_readdata,      --               .readdata
			rst       => rst_controller_reset_out_reset,                               --     reset_sink.reset
			blinky    => blinky_export                                                 --    conduit_end.export
		);

	iservo0 : component Computer_System_iServo0
		port map (
			clk        => system_pll_sys_clk_clk,                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_iservo0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_iservo0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_iservo0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_iservo0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_iservo0_s1_readdata,        --                    .readdata
			out_port   => iservo_control_0_export                       -- external_connection.export
		);

	iservo_0 : component Computer_System_iServo0
		port map (
			clk        => system_pll_sys_clk_clk,                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_iservo_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_iservo_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_iservo_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_iservo_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_iservo_0_s1_readdata,        --                    .readdata
			out_port   => iservo_control_1_export                        -- external_connection.export
		);

	video_lt24_controller_0 : component Computer_System_video_lt24_controller_0
		port map (
			clk           => video_pll_0_lcd_clk_clk,                                    --                clk.clk
			reset         => rst_controller_002_reset_out_reset,                         --              reset.reset
			ready         => video_pixel_buffer_dma_0_avalon_pixel_source_ready,         --   avalon_LT24_sink.ready
			startofpacket => video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket, --                   .startofpacket
			endofpacket   => video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket,   --                   .endofpacket
			data_in       => video_pixel_buffer_dma_0_avalon_pixel_source_data,          --                   .data
			data_in_valid => video_pixel_buffer_dma_0_avalon_pixel_source_valid,         --                   .valid
			lt24_lcd_on   => video_lt24_controller_0_lcd_on,                             -- external_interface.lcd_on
			lt24_reset_n  => video_lt24_controller_0_reset_n,                            --                   .reset_n
			csx           => video_lt24_controller_0_csx,                                --                   .csx
			data_to_lcd   => video_lt24_controller_0_data,                               --                   .data
			rdx           => video_lt24_controller_0_rdx,                                --                   .rdx
			wrx           => video_lt24_controller_0_wrx,                                --                   .wrx
			data_not_cmd  => video_lt24_controller_0_dcx                                 --                   .dcx
		);

	video_pixel_buffer_dma_0 : component Computer_System_video_pixel_buffer_dma_0
		port map (
			clk                  => video_pll_0_lcd_clk_clk,                                                    --                     clk.clk
			reset                => rst_controller_002_reset_out_reset,                                         --                   reset.reset
			master_readdatavalid => open,                                                                       -- avalon_pixel_dma_master.readdatavalid
			master_waitrequest   => open,                                                                       --                        .waitrequest
			master_address       => open,                                                                       --                        .address
			master_arbiterlock   => open,                                                                       --                        .lock
			master_read          => open,                                                                       --                        .read
			master_readdata      => open,                                                                       --                        .readdata
			slave_address        => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address,    --    avalon_control_slave.address
			slave_byteenable     => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable, --                        .byteenable
			slave_read           => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read,       --                        .read
			slave_write          => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write,      --                        .write
			slave_writedata      => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata,  --                        .writedata
			slave_readdata       => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata,   --                        .readdata
			stream_ready         => video_pixel_buffer_dma_0_avalon_pixel_source_ready,                         --     avalon_pixel_source.ready
			stream_startofpacket => video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket,                 --                        .startofpacket
			stream_endofpacket   => video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket,                   --                        .endofpacket
			stream_valid         => video_pixel_buffer_dma_0_avalon_pixel_source_valid,                         --                        .valid
			stream_data          => video_pixel_buffer_dma_0_avalon_pixel_source_data                           --                        .data
		);

	video_pll_0 : component Computer_System_video_pll_0
		port map (
			ref_clk_clk        => video_pll_0_ref_clk_clk,        --      ref_clk.clk
			ref_reset_reset    => video_pll_0_ref_reset_reset,    --    ref_reset.reset
			lcd_clk_clk        => video_pll_0_lcd_clk_clk,        --      lcd_clk.clk
			reset_source_reset => video_pll_0_reset_source_reset  -- reset_source.reset
		);

	nios2_custom_instruction_master_translator : component altera_customins_master_translator
		generic map (
			SHARED_COMB_AND_MULTI => 1
		)
		port map (
			ci_slave_dataa            => nios2_custom_instruction_master_dataa,                                --        ci_slave.dataa
			ci_slave_datab            => nios2_custom_instruction_master_datab,                                --                .datab
			ci_slave_result           => nios2_custom_instruction_master_result,                               --                .result
			ci_slave_n                => nios2_custom_instruction_master_n,                                    --                .n
			ci_slave_readra           => nios2_custom_instruction_master_readra,                               --                .readra
			ci_slave_readrb           => nios2_custom_instruction_master_readrb,                               --                .readrb
			ci_slave_writerc          => nios2_custom_instruction_master_writerc,                              --                .writerc
			ci_slave_a                => nios2_custom_instruction_master_a,                                    --                .a
			ci_slave_b                => nios2_custom_instruction_master_b,                                    --                .b
			ci_slave_c                => nios2_custom_instruction_master_c,                                    --                .c
			ci_slave_ipending         => nios2_custom_instruction_master_ipending,                             --                .ipending
			ci_slave_estatus          => nios2_custom_instruction_master_estatus,                              --                .estatus
			ci_slave_multi_clk        => nios2_custom_instruction_master_clk,                                  --                .clk
			ci_slave_multi_reset      => nios2_custom_instruction_master_reset,                                --                .reset
			ci_slave_multi_clken      => nios2_custom_instruction_master_clk_en,                               --                .clk_en
			ci_slave_multi_reset_req  => nios2_custom_instruction_master_reset_req,                            --                .reset_req
			ci_slave_multi_start      => nios2_custom_instruction_master_start,                                --                .start
			ci_slave_multi_done       => nios2_custom_instruction_master_done,                                 --                .done
			comb_ci_master_dataa      => open,                                                                 --  comb_ci_master.dataa
			comb_ci_master_datab      => open,                                                                 --                .datab
			comb_ci_master_result     => open,                                                                 --                .result
			comb_ci_master_n          => open,                                                                 --                .n
			comb_ci_master_readra     => open,                                                                 --                .readra
			comb_ci_master_readrb     => open,                                                                 --                .readrb
			comb_ci_master_writerc    => open,                                                                 --                .writerc
			comb_ci_master_a          => open,                                                                 --                .a
			comb_ci_master_b          => open,                                                                 --                .b
			comb_ci_master_c          => open,                                                                 --                .c
			comb_ci_master_ipending   => open,                                                                 --                .ipending
			comb_ci_master_estatus    => open,                                                                 --                .estatus
			multi_ci_master_clk       => nios2_custom_instruction_master_translator_multi_ci_master_clk,       -- multi_ci_master.clk
			multi_ci_master_reset     => nios2_custom_instruction_master_translator_multi_ci_master_reset,     --                .reset
			multi_ci_master_clken     => nios2_custom_instruction_master_translator_multi_ci_master_clk_en,    --                .clk_en
			multi_ci_master_reset_req => nios2_custom_instruction_master_translator_multi_ci_master_reset_req, --                .reset_req
			multi_ci_master_start     => nios2_custom_instruction_master_translator_multi_ci_master_start,     --                .start
			multi_ci_master_done      => nios2_custom_instruction_master_translator_multi_ci_master_done,      --                .done
			multi_ci_master_dataa     => nios2_custom_instruction_master_translator_multi_ci_master_dataa,     --                .dataa
			multi_ci_master_datab     => nios2_custom_instruction_master_translator_multi_ci_master_datab,     --                .datab
			multi_ci_master_result    => nios2_custom_instruction_master_translator_multi_ci_master_result,    --                .result
			multi_ci_master_n         => nios2_custom_instruction_master_translator_multi_ci_master_n,         --                .n
			multi_ci_master_readra    => nios2_custom_instruction_master_translator_multi_ci_master_readra,    --                .readra
			multi_ci_master_readrb    => nios2_custom_instruction_master_translator_multi_ci_master_readrb,    --                .readrb
			multi_ci_master_writerc   => nios2_custom_instruction_master_translator_multi_ci_master_writerc,   --                .writerc
			multi_ci_master_a         => nios2_custom_instruction_master_translator_multi_ci_master_a,         --                .a
			multi_ci_master_b         => nios2_custom_instruction_master_translator_multi_ci_master_b,         --                .b
			multi_ci_master_c         => nios2_custom_instruction_master_translator_multi_ci_master_c,         --                .c
			ci_slave_multi_dataa      => "00000000000000000000000000000000",                                   --     (terminated)
			ci_slave_multi_datab      => "00000000000000000000000000000000",                                   --     (terminated)
			ci_slave_multi_result     => open,                                                                 --     (terminated)
			ci_slave_multi_n          => "00000000",                                                           --     (terminated)
			ci_slave_multi_readra     => '0',                                                                  --     (terminated)
			ci_slave_multi_readrb     => '0',                                                                  --     (terminated)
			ci_slave_multi_writerc    => '0',                                                                  --     (terminated)
			ci_slave_multi_a          => "00000",                                                              --     (terminated)
			ci_slave_multi_b          => "00000",                                                              --     (terminated)
			ci_slave_multi_c          => "00000"                                                               --     (terminated)
		);

	nios2_custom_instruction_master_multi_xconnect : component Computer_System_Nios2_custom_instruction_master_multi_xconnect
		port map (
			ci_slave_dataa       => nios2_custom_instruction_master_translator_multi_ci_master_dataa,     --   ci_slave.dataa
			ci_slave_datab       => nios2_custom_instruction_master_translator_multi_ci_master_datab,     --           .datab
			ci_slave_result      => nios2_custom_instruction_master_translator_multi_ci_master_result,    --           .result
			ci_slave_n           => nios2_custom_instruction_master_translator_multi_ci_master_n,         --           .n
			ci_slave_readra      => nios2_custom_instruction_master_translator_multi_ci_master_readra,    --           .readra
			ci_slave_readrb      => nios2_custom_instruction_master_translator_multi_ci_master_readrb,    --           .readrb
			ci_slave_writerc     => nios2_custom_instruction_master_translator_multi_ci_master_writerc,   --           .writerc
			ci_slave_a           => nios2_custom_instruction_master_translator_multi_ci_master_a,         --           .a
			ci_slave_b           => nios2_custom_instruction_master_translator_multi_ci_master_b,         --           .b
			ci_slave_c           => nios2_custom_instruction_master_translator_multi_ci_master_c,         --           .c
			ci_slave_ipending    => open,                                                                 --           .ipending
			ci_slave_estatus     => open,                                                                 --           .estatus
			ci_slave_clk         => nios2_custom_instruction_master_translator_multi_ci_master_clk,       --           .clk
			ci_slave_reset       => nios2_custom_instruction_master_translator_multi_ci_master_reset,     --           .reset
			ci_slave_clken       => nios2_custom_instruction_master_translator_multi_ci_master_clk_en,    --           .clk_en
			ci_slave_reset_req   => nios2_custom_instruction_master_translator_multi_ci_master_reset_req, --           .reset_req
			ci_slave_start       => nios2_custom_instruction_master_translator_multi_ci_master_start,     --           .start
			ci_slave_done        => nios2_custom_instruction_master_translator_multi_ci_master_done,      --           .done
			ci_master0_dataa     => nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa,      -- ci_master0.dataa
			ci_master0_datab     => nios2_custom_instruction_master_multi_xconnect_ci_master0_datab,      --           .datab
			ci_master0_result    => nios2_custom_instruction_master_multi_xconnect_ci_master0_result,     --           .result
			ci_master0_n         => nios2_custom_instruction_master_multi_xconnect_ci_master0_n,          --           .n
			ci_master0_readra    => nios2_custom_instruction_master_multi_xconnect_ci_master0_readra,     --           .readra
			ci_master0_readrb    => nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb,     --           .readrb
			ci_master0_writerc   => nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc,    --           .writerc
			ci_master0_a         => nios2_custom_instruction_master_multi_xconnect_ci_master0_a,          --           .a
			ci_master0_b         => nios2_custom_instruction_master_multi_xconnect_ci_master0_b,          --           .b
			ci_master0_c         => nios2_custom_instruction_master_multi_xconnect_ci_master0_c,          --           .c
			ci_master0_ipending  => nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending,   --           .ipending
			ci_master0_estatus   => nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus,    --           .estatus
			ci_master0_clk       => nios2_custom_instruction_master_multi_xconnect_ci_master0_clk,        --           .clk
			ci_master0_reset     => nios2_custom_instruction_master_multi_xconnect_ci_master0_reset,      --           .reset
			ci_master0_clken     => nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en,     --           .clk_en
			ci_master0_reset_req => nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req,  --           .reset_req
			ci_master0_start     => nios2_custom_instruction_master_multi_xconnect_ci_master0_start,      --           .start
			ci_master0_done      => nios2_custom_instruction_master_multi_xconnect_ci_master0_done        --           .done
		);

	nios2_custom_instruction_master_multi_slave_translator0 : component altera_customins_slave_translator
		generic map (
			N_WIDTH          => 2,
			USE_DONE         => 1,
			NUM_FIXED_CYCLES => 1
		)
		port map (
			ci_slave_dataa      => nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa,          --  ci_slave.dataa
			ci_slave_datab      => nios2_custom_instruction_master_multi_xconnect_ci_master0_datab,          --          .datab
			ci_slave_result     => nios2_custom_instruction_master_multi_xconnect_ci_master0_result,         --          .result
			ci_slave_n          => nios2_custom_instruction_master_multi_xconnect_ci_master0_n,              --          .n
			ci_slave_readra     => nios2_custom_instruction_master_multi_xconnect_ci_master0_readra,         --          .readra
			ci_slave_readrb     => nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb,         --          .readrb
			ci_slave_writerc    => nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc,        --          .writerc
			ci_slave_a          => nios2_custom_instruction_master_multi_xconnect_ci_master0_a,              --          .a
			ci_slave_b          => nios2_custom_instruction_master_multi_xconnect_ci_master0_b,              --          .b
			ci_slave_c          => nios2_custom_instruction_master_multi_xconnect_ci_master0_c,              --          .c
			ci_slave_ipending   => nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending,       --          .ipending
			ci_slave_estatus    => nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus,        --          .estatus
			ci_slave_clk        => nios2_custom_instruction_master_multi_xconnect_ci_master0_clk,            --          .clk
			ci_slave_clken      => nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en,         --          .clk_en
			ci_slave_reset_req  => nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req,      --          .reset_req
			ci_slave_reset      => nios2_custom_instruction_master_multi_xconnect_ci_master0_reset,          --          .reset
			ci_slave_start      => nios2_custom_instruction_master_multi_xconnect_ci_master0_start,          --          .start
			ci_slave_done       => nios2_custom_instruction_master_multi_xconnect_ci_master0_done,           --          .done
			ci_master_dataa     => nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa,  -- ci_master.dataa
			ci_master_datab     => nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab,  --          .datab
			ci_master_result    => nios2_custom_instruction_master_multi_slave_translator0_ci_master_result, --          .result
			ci_master_n         => nios2_custom_instruction_master_multi_slave_translator0_ci_master_n,      --          .n
			ci_master_clk       => nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk,    --          .clk
			ci_master_clken     => nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en, --          .clk_en
			ci_master_reset     => nios2_custom_instruction_master_multi_slave_translator0_ci_master_reset,  --          .reset
			ci_master_start     => nios2_custom_instruction_master_multi_slave_translator0_ci_master_start,  --          .start
			ci_master_done      => nios2_custom_instruction_master_multi_slave_translator0_ci_master_done,   --          .done
			ci_master_readra    => open,                                                                     -- (terminated)
			ci_master_readrb    => open,                                                                     -- (terminated)
			ci_master_writerc   => open,                                                                     -- (terminated)
			ci_master_a         => open,                                                                     -- (terminated)
			ci_master_b         => open,                                                                     -- (terminated)
			ci_master_c         => open,                                                                     -- (terminated)
			ci_master_ipending  => open,                                                                     -- (terminated)
			ci_master_estatus   => open,                                                                     -- (terminated)
			ci_master_reset_req => open                                                                      -- (terminated)
		);

	mm_interconnect_0 : component Computer_System_mm_interconnect_0
		port map (
			System_PLL_sys_clk_clk                                     => system_pll_sys_clk_clk,                                                     --                                   System_PLL_sys_clk.clk
			video_pll_0_lcd_clk_clk                                    => video_pll_0_lcd_clk_clk,                                                    --                                  video_pll_0_lcd_clk.clk
			ADC_reset_reset_bridge_in_reset_reset                      => rst_controller_reset_out_reset,                                             --                      ADC_reset_reset_bridge_in_reset.reset
			JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset  => rst_controller_reset_out_reset,                                             --  JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset.reset
			Nios2_reset_reset_bridge_in_reset_reset                    => rst_controller_001_reset_out_reset,                                         --                    Nios2_reset_reset_bridge_in_reset.reset
			video_pixel_buffer_dma_0_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                                         -- video_pixel_buffer_dma_0_reset_reset_bridge_in_reset.reset
			JTAG_to_FPGA_Bridge_master_address                         => jtag_to_fpga_bridge_master_address,                                         --                           JTAG_to_FPGA_Bridge_master.address
			JTAG_to_FPGA_Bridge_master_waitrequest                     => jtag_to_fpga_bridge_master_waitrequest,                                     --                                                     .waitrequest
			JTAG_to_FPGA_Bridge_master_byteenable                      => jtag_to_fpga_bridge_master_byteenable,                                      --                                                     .byteenable
			JTAG_to_FPGA_Bridge_master_read                            => jtag_to_fpga_bridge_master_read,                                            --                                                     .read
			JTAG_to_FPGA_Bridge_master_readdata                        => jtag_to_fpga_bridge_master_readdata,                                        --                                                     .readdata
			JTAG_to_FPGA_Bridge_master_readdatavalid                   => jtag_to_fpga_bridge_master_readdatavalid,                                   --                                                     .readdatavalid
			JTAG_to_FPGA_Bridge_master_write                           => jtag_to_fpga_bridge_master_write,                                           --                                                     .write
			JTAG_to_FPGA_Bridge_master_writedata                       => jtag_to_fpga_bridge_master_writedata,                                       --                                                     .writedata
			Nios2_data_master_address                                  => nios2_data_master_address,                                                  --                                    Nios2_data_master.address
			Nios2_data_master_waitrequest                              => nios2_data_master_waitrequest,                                              --                                                     .waitrequest
			Nios2_data_master_byteenable                               => nios2_data_master_byteenable,                                               --                                                     .byteenable
			Nios2_data_master_read                                     => nios2_data_master_read,                                                     --                                                     .read
			Nios2_data_master_readdata                                 => nios2_data_master_readdata,                                                 --                                                     .readdata
			Nios2_data_master_write                                    => nios2_data_master_write,                                                    --                                                     .write
			Nios2_data_master_writedata                                => nios2_data_master_writedata,                                                --                                                     .writedata
			Nios2_data_master_debugaccess                              => nios2_data_master_debugaccess,                                              --                                                     .debugaccess
			Nios2_instruction_master_address                           => nios2_instruction_master_address,                                           --                             Nios2_instruction_master.address
			Nios2_instruction_master_waitrequest                       => nios2_instruction_master_waitrequest,                                       --                                                     .waitrequest
			Nios2_instruction_master_read                              => nios2_instruction_master_read,                                              --                                                     .read
			Nios2_instruction_master_readdata                          => nios2_instruction_master_readdata,                                          --                                                     .readdata
			ADC_adc_slave_address                                      => mm_interconnect_0_adc_adc_slave_address,                                    --                                        ADC_adc_slave.address
			ADC_adc_slave_write                                        => mm_interconnect_0_adc_adc_slave_write,                                      --                                                     .write
			ADC_adc_slave_read                                         => mm_interconnect_0_adc_adc_slave_read,                                       --                                                     .read
			ADC_adc_slave_readdata                                     => mm_interconnect_0_adc_adc_slave_readdata,                                   --                                                     .readdata
			ADC_adc_slave_writedata                                    => mm_interconnect_0_adc_adc_slave_writedata,                                  --                                                     .writedata
			ADC_adc_slave_waitrequest                                  => mm_interconnect_0_adc_adc_slave_waitrequest,                                --                                                     .waitrequest
			Arduino_GPIO_s1_address                                    => mm_interconnect_0_arduino_gpio_s1_address,                                  --                                      Arduino_GPIO_s1.address
			Arduino_GPIO_s1_write                                      => mm_interconnect_0_arduino_gpio_s1_write,                                    --                                                     .write
			Arduino_GPIO_s1_readdata                                   => mm_interconnect_0_arduino_gpio_s1_readdata,                                 --                                                     .readdata
			Arduino_GPIO_s1_writedata                                  => mm_interconnect_0_arduino_gpio_s1_writedata,                                --                                                     .writedata
			Arduino_GPIO_s1_chipselect                                 => mm_interconnect_0_arduino_gpio_s1_chipselect,                               --                                                     .chipselect
			Arduino_Reset_N_s1_address                                 => mm_interconnect_0_arduino_reset_n_s1_address,                               --                                   Arduino_Reset_N_s1.address
			Arduino_Reset_N_s1_write                                   => mm_interconnect_0_arduino_reset_n_s1_write,                                 --                                                     .write
			Arduino_Reset_N_s1_readdata                                => mm_interconnect_0_arduino_reset_n_s1_readdata,                              --                                                     .readdata
			Arduino_Reset_N_s1_writedata                               => mm_interconnect_0_arduino_reset_n_s1_writedata,                             --                                                     .writedata
			Arduino_Reset_N_s1_chipselect                              => mm_interconnect_0_arduino_reset_n_s1_chipselect,                            --                                                     .chipselect
			blinky_test_0_avalon_slave_0_address                       => mm_interconnect_0_blinky_test_0_avalon_slave_0_address,                     --                         blinky_test_0_avalon_slave_0.address
			blinky_test_0_avalon_slave_0_write                         => mm_interconnect_0_blinky_test_0_avalon_slave_0_write,                       --                                                     .write
			blinky_test_0_avalon_slave_0_read                          => mm_interconnect_0_blinky_test_0_avalon_slave_0_read,                        --                                                     .read
			blinky_test_0_avalon_slave_0_readdata                      => mm_interconnect_0_blinky_test_0_avalon_slave_0_readdata,                    --                                                     .readdata
			blinky_test_0_avalon_slave_0_writedata                     => mm_interconnect_0_blinky_test_0_avalon_slave_0_writedata,                   --                                                     .writedata
			blinky_test_0_avalon_slave_0_byteenable                    => mm_interconnect_0_blinky_test_0_avalon_slave_0_byteenable,                  --                                                     .byteenable
			Expansion_JP1_s1_address                                   => mm_interconnect_0_expansion_jp1_s1_address,                                 --                                     Expansion_JP1_s1.address
			Expansion_JP1_s1_write                                     => mm_interconnect_0_expansion_jp1_s1_write,                                   --                                                     .write
			Expansion_JP1_s1_readdata                                  => mm_interconnect_0_expansion_jp1_s1_readdata,                                --                                                     .readdata
			Expansion_JP1_s1_writedata                                 => mm_interconnect_0_expansion_jp1_s1_writedata,                               --                                                     .writedata
			Expansion_JP1_s1_chipselect                                => mm_interconnect_0_expansion_jp1_s1_chipselect,                              --                                                     .chipselect
			HEX3_HEX0_s1_address                                       => mm_interconnect_0_hex3_hex0_s1_address,                                     --                                         HEX3_HEX0_s1.address
			HEX3_HEX0_s1_write                                         => mm_interconnect_0_hex3_hex0_s1_write,                                       --                                                     .write
			HEX3_HEX0_s1_readdata                                      => mm_interconnect_0_hex3_hex0_s1_readdata,                                    --                                                     .readdata
			HEX3_HEX0_s1_writedata                                     => mm_interconnect_0_hex3_hex0_s1_writedata,                                   --                                                     .writedata
			HEX3_HEX0_s1_chipselect                                    => mm_interconnect_0_hex3_hex0_s1_chipselect,                                  --                                                     .chipselect
			HEX5_HEX4_s1_address                                       => mm_interconnect_0_hex5_hex4_s1_address,                                     --                                         HEX5_HEX4_s1.address
			HEX5_HEX4_s1_write                                         => mm_interconnect_0_hex5_hex4_s1_write,                                       --                                                     .write
			HEX5_HEX4_s1_readdata                                      => mm_interconnect_0_hex5_hex4_s1_readdata,                                    --                                                     .readdata
			HEX5_HEX4_s1_writedata                                     => mm_interconnect_0_hex5_hex4_s1_writedata,                                   --                                                     .writedata
			HEX5_HEX4_s1_chipselect                                    => mm_interconnect_0_hex5_hex4_s1_chipselect,                                  --                                                     .chipselect
			Interval_Timer_s1_address                                  => mm_interconnect_0_interval_timer_s1_address,                                --                                    Interval_Timer_s1.address
			Interval_Timer_s1_write                                    => mm_interconnect_0_interval_timer_s1_write,                                  --                                                     .write
			Interval_Timer_s1_readdata                                 => mm_interconnect_0_interval_timer_s1_readdata,                               --                                                     .readdata
			Interval_Timer_s1_writedata                                => mm_interconnect_0_interval_timer_s1_writedata,                              --                                                     .writedata
			Interval_Timer_s1_chipselect                               => mm_interconnect_0_interval_timer_s1_chipselect,                             --                                                     .chipselect
			Interval_Timer_2_s1_address                                => mm_interconnect_0_interval_timer_2_s1_address,                              --                                  Interval_Timer_2_s1.address
			Interval_Timer_2_s1_write                                  => mm_interconnect_0_interval_timer_2_s1_write,                                --                                                     .write
			Interval_Timer_2_s1_readdata                               => mm_interconnect_0_interval_timer_2_s1_readdata,                             --                                                     .readdata
			Interval_Timer_2_s1_writedata                              => mm_interconnect_0_interval_timer_2_s1_writedata,                            --                                                     .writedata
			Interval_Timer_2_s1_chipselect                             => mm_interconnect_0_interval_timer_2_s1_chipselect,                           --                                                     .chipselect
			iServo0_s1_address                                         => mm_interconnect_0_iservo0_s1_address,                                       --                                           iServo0_s1.address
			iServo0_s1_write                                           => mm_interconnect_0_iservo0_s1_write,                                         --                                                     .write
			iServo0_s1_readdata                                        => mm_interconnect_0_iservo0_s1_readdata,                                      --                                                     .readdata
			iServo0_s1_writedata                                       => mm_interconnect_0_iservo0_s1_writedata,                                     --                                                     .writedata
			iServo0_s1_chipselect                                      => mm_interconnect_0_iservo0_s1_chipselect,                                    --                                                     .chipselect
			iServo_0_s1_address                                        => mm_interconnect_0_iservo_0_s1_address,                                      --                                          iServo_0_s1.address
			iServo_0_s1_write                                          => mm_interconnect_0_iservo_0_s1_write,                                        --                                                     .write
			iServo_0_s1_readdata                                       => mm_interconnect_0_iservo_0_s1_readdata,                                     --                                                     .readdata
			iServo_0_s1_writedata                                      => mm_interconnect_0_iservo_0_s1_writedata,                                    --                                                     .writedata
			iServo_0_s1_chipselect                                     => mm_interconnect_0_iservo_0_s1_chipselect,                                   --                                                     .chipselect
			JTAG_UART_avalon_jtag_slave_address                        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,                      --                          JTAG_UART_avalon_jtag_slave.address
			JTAG_UART_avalon_jtag_slave_write                          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,                        --                                                     .write
			JTAG_UART_avalon_jtag_slave_read                           => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,                         --                                                     .read
			JTAG_UART_avalon_jtag_slave_readdata                       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,                     --                                                     .readdata
			JTAG_UART_avalon_jtag_slave_writedata                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,                    --                                                     .writedata
			JTAG_UART_avalon_jtag_slave_waitrequest                    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,                  --                                                     .waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,                   --                                                     .chipselect
			LEDs_s1_address                                            => mm_interconnect_0_leds_s1_address,                                          --                                              LEDs_s1.address
			LEDs_s1_write                                              => mm_interconnect_0_leds_s1_write,                                            --                                                     .write
			LEDs_s1_readdata                                           => mm_interconnect_0_leds_s1_readdata,                                         --                                                     .readdata
			LEDs_s1_writedata                                          => mm_interconnect_0_leds_s1_writedata,                                        --                                                     .writedata
			LEDs_s1_chipselect                                         => mm_interconnect_0_leds_s1_chipselect,                                       --                                                     .chipselect
			Nios2_debug_mem_slave_address                              => mm_interconnect_0_nios2_debug_mem_slave_address,                            --                                Nios2_debug_mem_slave.address
			Nios2_debug_mem_slave_write                                => mm_interconnect_0_nios2_debug_mem_slave_write,                              --                                                     .write
			Nios2_debug_mem_slave_read                                 => mm_interconnect_0_nios2_debug_mem_slave_read,                               --                                                     .read
			Nios2_debug_mem_slave_readdata                             => mm_interconnect_0_nios2_debug_mem_slave_readdata,                           --                                                     .readdata
			Nios2_debug_mem_slave_writedata                            => mm_interconnect_0_nios2_debug_mem_slave_writedata,                          --                                                     .writedata
			Nios2_debug_mem_slave_byteenable                           => mm_interconnect_0_nios2_debug_mem_slave_byteenable,                         --                                                     .byteenable
			Nios2_debug_mem_slave_waitrequest                          => mm_interconnect_0_nios2_debug_mem_slave_waitrequest,                        --                                                     .waitrequest
			Nios2_debug_mem_slave_debugaccess                          => mm_interconnect_0_nios2_debug_mem_slave_debugaccess,                        --                                                     .debugaccess
			Onchip_SRAM_s1_address                                     => mm_interconnect_0_onchip_sram_s1_address,                                   --                                       Onchip_SRAM_s1.address
			Onchip_SRAM_s1_write                                       => mm_interconnect_0_onchip_sram_s1_write,                                     --                                                     .write
			Onchip_SRAM_s1_readdata                                    => mm_interconnect_0_onchip_sram_s1_readdata,                                  --                                                     .readdata
			Onchip_SRAM_s1_writedata                                   => mm_interconnect_0_onchip_sram_s1_writedata,                                 --                                                     .writedata
			Onchip_SRAM_s1_byteenable                                  => mm_interconnect_0_onchip_sram_s1_byteenable,                                --                                                     .byteenable
			Onchip_SRAM_s1_chipselect                                  => mm_interconnect_0_onchip_sram_s1_chipselect,                                --                                                     .chipselect
			Onchip_SRAM_s1_clken                                       => mm_interconnect_0_onchip_sram_s1_clken,                                     --                                                     .clken
			Onchip_SRAM_s2_address                                     => mm_interconnect_0_onchip_sram_s2_address,                                   --                                       Onchip_SRAM_s2.address
			Onchip_SRAM_s2_write                                       => mm_interconnect_0_onchip_sram_s2_write,                                     --                                                     .write
			Onchip_SRAM_s2_readdata                                    => mm_interconnect_0_onchip_sram_s2_readdata,                                  --                                                     .readdata
			Onchip_SRAM_s2_writedata                                   => mm_interconnect_0_onchip_sram_s2_writedata,                                 --                                                     .writedata
			Onchip_SRAM_s2_byteenable                                  => mm_interconnect_0_onchip_sram_s2_byteenable,                                --                                                     .byteenable
			Onchip_SRAM_s2_chipselect                                  => mm_interconnect_0_onchip_sram_s2_chipselect,                                --                                                     .chipselect
			Onchip_SRAM_s2_clken                                       => mm_interconnect_0_onchip_sram_s2_clken,                                     --                                                     .clken
			Pushbuttons_s1_address                                     => mm_interconnect_0_pushbuttons_s1_address,                                   --                                       Pushbuttons_s1.address
			Pushbuttons_s1_write                                       => mm_interconnect_0_pushbuttons_s1_write,                                     --                                                     .write
			Pushbuttons_s1_readdata                                    => mm_interconnect_0_pushbuttons_s1_readdata,                                  --                                                     .readdata
			Pushbuttons_s1_writedata                                   => mm_interconnect_0_pushbuttons_s1_writedata,                                 --                                                     .writedata
			Pushbuttons_s1_chipselect                                  => mm_interconnect_0_pushbuttons_s1_chipselect,                                --                                                     .chipselect
			SDRAM_s1_address                                           => mm_interconnect_0_sdram_s1_address,                                         --                                             SDRAM_s1.address
			SDRAM_s1_write                                             => mm_interconnect_0_sdram_s1_write,                                           --                                                     .write
			SDRAM_s1_read                                              => mm_interconnect_0_sdram_s1_read,                                            --                                                     .read
			SDRAM_s1_readdata                                          => mm_interconnect_0_sdram_s1_readdata,                                        --                                                     .readdata
			SDRAM_s1_writedata                                         => mm_interconnect_0_sdram_s1_writedata,                                       --                                                     .writedata
			SDRAM_s1_byteenable                                        => mm_interconnect_0_sdram_s1_byteenable,                                      --                                                     .byteenable
			SDRAM_s1_readdatavalid                                     => mm_interconnect_0_sdram_s1_readdatavalid,                                   --                                                     .readdatavalid
			SDRAM_s1_waitrequest                                       => mm_interconnect_0_sdram_s1_waitrequest,                                     --                                                     .waitrequest
			SDRAM_s1_chipselect                                        => mm_interconnect_0_sdram_s1_chipselect,                                      --                                                     .chipselect
			Servo0_servo_control_slave_address                         => mm_interconnect_0_servo0_servo_control_slave_address,                       --                           Servo0_servo_control_slave.address
			Servo0_servo_control_slave_write                           => mm_interconnect_0_servo0_servo_control_slave_write,                         --                                                     .write
			Servo0_servo_control_slave_read                            => mm_interconnect_0_servo0_servo_control_slave_read,                          --                                                     .read
			Servo0_servo_control_slave_readdata                        => mm_interconnect_0_servo0_servo_control_slave_readdata,                      --                                                     .readdata
			Servo0_servo_control_slave_writedata                       => mm_interconnect_0_servo0_servo_control_slave_writedata,                     --                                                     .writedata
			Servo0_servo_control_slave_byteenable                      => mm_interconnect_0_servo0_servo_control_slave_byteenable,                    --                                                     .byteenable
			Servo1_servo_control_slave_address                         => mm_interconnect_0_servo1_servo_control_slave_address,                       --                           Servo1_servo_control_slave.address
			Servo1_servo_control_slave_write                           => mm_interconnect_0_servo1_servo_control_slave_write,                         --                                                     .write
			Servo1_servo_control_slave_read                            => mm_interconnect_0_servo1_servo_control_slave_read,                          --                                                     .read
			Servo1_servo_control_slave_readdata                        => mm_interconnect_0_servo1_servo_control_slave_readdata,                      --                                                     .readdata
			Servo1_servo_control_slave_writedata                       => mm_interconnect_0_servo1_servo_control_slave_writedata,                     --                                                     .writedata
			Servo1_servo_control_slave_byteenable                      => mm_interconnect_0_servo1_servo_control_slave_byteenable,                    --                                                     .byteenable
			Slider_Switches_s1_address                                 => mm_interconnect_0_slider_switches_s1_address,                               --                                   Slider_Switches_s1.address
			Slider_Switches_s1_readdata                                => mm_interconnect_0_slider_switches_s1_readdata,                              --                                                     .readdata
			SysID_control_slave_address                                => mm_interconnect_0_sysid_control_slave_address,                              --                                  SysID_control_slave.address
			SysID_control_slave_readdata                               => mm_interconnect_0_sysid_control_slave_readdata,                             --                                                     .readdata
			video_pixel_buffer_dma_0_avalon_control_slave_address      => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address,    --        video_pixel_buffer_dma_0_avalon_control_slave.address
			video_pixel_buffer_dma_0_avalon_control_slave_write        => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write,      --                                                     .write
			video_pixel_buffer_dma_0_avalon_control_slave_read         => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read,       --                                                     .read
			video_pixel_buffer_dma_0_avalon_control_slave_readdata     => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata,   --                                                     .readdata
			video_pixel_buffer_dma_0_avalon_control_slave_writedata    => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata,  --                                                     .writedata
			video_pixel_buffer_dma_0_avalon_control_slave_byteenable   => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable  --                                                     .byteenable
		);

	irq_mapper : component Computer_System_irq_mapper
		port map (
			clk           => system_pll_sys_clk_clk,             --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,           -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,           -- receiver5.irq
			sender_irq    => nios2_irq_irq                       --    sender.irq
		);

	rst_controller : component computer_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => system_pll_reset_source_reset,      -- reset_in0.reset
			clk            => system_pll_sys_clk_clk,             --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component computer_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_debug_reset_request_reset,    -- reset_in0.reset
			reset_in1      => system_pll_reset_source_reset,      -- reset_in1.reset
			clk            => system_pll_sys_clk_clk,             --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component computer_system_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => video_pll_0_reset_source_reset,     -- reset_in0.reset
			clk            => video_pll_0_lcd_clk_clk,            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_leds_s1_write_ports_inv <= not mm_interconnect_0_leds_s1_write;

	mm_interconnect_0_hex3_hex0_s1_write_ports_inv <= not mm_interconnect_0_hex3_hex0_s1_write;

	mm_interconnect_0_hex5_hex4_s1_write_ports_inv <= not mm_interconnect_0_hex5_hex4_s1_write;

	mm_interconnect_0_pushbuttons_s1_write_ports_inv <= not mm_interconnect_0_pushbuttons_s1_write;

	mm_interconnect_0_expansion_jp1_s1_write_ports_inv <= not mm_interconnect_0_expansion_jp1_s1_write;

	mm_interconnect_0_arduino_gpio_s1_write_ports_inv <= not mm_interconnect_0_arduino_gpio_s1_write;

	mm_interconnect_0_arduino_reset_n_s1_write_ports_inv <= not mm_interconnect_0_arduino_reset_n_s1_write;

	mm_interconnect_0_interval_timer_s1_write_ports_inv <= not mm_interconnect_0_interval_timer_s1_write;

	mm_interconnect_0_interval_timer_2_s1_write_ports_inv <= not mm_interconnect_0_interval_timer_2_s1_write;

	mm_interconnect_0_iservo0_s1_write_ports_inv <= not mm_interconnect_0_iservo0_s1_write;

	mm_interconnect_0_iservo_0_s1_write_ports_inv <= not mm_interconnect_0_iservo_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of Computer_System
